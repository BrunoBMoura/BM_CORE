/*
clk_write - clock
clk_read - auto clock
proc_num - 0 or 1, indicates if it's the OS or one of the processes that's beeing executed
write_flag - flag for data storage
write_os - only using during BIOS operations, write flag for OS instructions
input_data - data to be stored
write_address - self explanatory
read_address - self explanatory
instr_mem_out - output value of InstrMem
*/

module Instruction_memory
#(
	parameter DATA_WIDTH = 32, 
	parameter REGION_WIDTH = 11
)
(
	input clk_write, clk_read, proc_num, write_flag, write_os,
	input [(DATA_WIDTH-1):0] write_address, read_address,
	input [(DATA_WIDTH-1):0] input_data,
	output [(DATA_WIDTH-1):0] instr_mem_out
);
	
	reg [(DATA_WIDTH-1):0] proc_mem[(2**REGION_WIDTH-1):0];
	reg [(DATA_WIDTH-1):0] os_mem[(2**REGION_WIDTH-1):0];
	reg [(DATA_WIDTH-1):0] data_os_out, data_proc_out;
  
	always @ ( posedge clk_write ) 
	begin
		if( write_flag )
		begin
			if( write_os ) 
				os_mem[ write_address ] <= input_data;
			else
				proc_mem[ write_address ] <= input_data;
		end
			
	end
	
	always @ ( posedge clk_read )
	begin
		data_os_out <= os_mem[ read_address ];
		data_proc_out <= proc_mem[ read_address ];
	end

	assign instr_mem_out = (proc_num == 1'b0) ? data_os_out : data_proc_out;
	
 endmodule 
 
		
	
		/*
		instrmem[0] <= 32'b010000_00000_11110_0000000000000000; // $sp = 0
		instrmem[1] <= 32'b010100_00000000000000000100010110; // jump to 278(main)
		instrmem[2] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[3] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[4] <= 32'b010001_00000_00001_0000000000000010; // m[r[0] + 2] = r[1]
		instrmem[5] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[6] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[7] <= 32'b010001_00000_00001_0000000000000001; // m[r[0] + 1] = r[1]
		instrmem[8] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[9] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[10] <= 32'b010001_00000_00001_0000000000000000; // m[r[0] + 0] = r[1]
		instrmem[11] <= 32'b001111_00000_00001_0000000000000001; // r[1] = m[r[0] + 1]
		instrmem[12] <= 32'b010001_00000_00001_0000000000000101; // m[r[0] + 5] = r[1]
		instrmem[13] <= 32'b001111_00000_00001_0000000000000000; // r[1] = m[r[0] + 0]
		instrmem[14] <= 32'b001111_00000_00010_0000000000000001; // r[2] = m[r[0] + 1]
		instrmem[15] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		instrmem[16] <= 32'b001111_00001_00010_0000000000000000; // r[2] = m[r[1] + 0]
		instrmem[17] <= 32'b010001_00000_00010_0000000000000100; // m[r[0] + 4] = r[2]
		instrmem[18] <= 32'b001111_00000_00001_0000000000000001; // r[1] = m[r[0] + 1]
		instrmem[19] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		instrmem[20] <= 32'b010001_00000_00001_0000000000000011; // m[r[0] + 3] = r[1]
		instrmem[21] <= 32'b001111_00000_00001_0000000000000011; // r[1] = m[r[0] + 3]
		instrmem[22] <= 32'b001111_00000_00010_0000000000000010; // r[2] = m[r[0] + 2]
		instrmem[23] <= 32'b000110_00001_00010_00011_00000_000000; // (r[1] < r[2]) ? r[3] = 1 : r[3] = 0
		instrmem[24] <= 32'b010010_00000_00011_0000000000101011; // if(r[0] == r[3]) jump to 43(L3)
		instrmem[25] <= 32'b001111_00000_00001_0000000000000000; // r[1] = m[r[0] + 0]
		instrmem[26] <= 32'b001111_00000_00010_0000000000000011; // r[2] = m[r[0] + 3]
		instrmem[27] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		instrmem[28] <= 32'b001111_00001_00010_0000000000000000; // r[2] = m[r[1] + 0]
		instrmem[29] <= 32'b001111_00000_00001_0000000000000100; // r[1] = m[r[0] + 4]
		instrmem[30] <= 32'b000110_00010_00001_00100_00000_000000; // (r[2] < r[1]) ? r[4] = 1 : r[4] = 0
		instrmem[31] <= 32'b010010_00000_00100_0000000000100111; // if(r[0] == r[4]) jump to 39(L5)
		instrmem[32] <= 32'b001111_00000_00001_0000000000000000; // r[1] = m[r[0] + 0]
		instrmem[33] <= 32'b001111_00000_00010_0000000000000011; // r[2] = m[r[0] + 3]
		instrmem[34] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		instrmem[35] <= 32'b001111_00001_00010_0000000000000000; // r[2] = m[r[1] + 0]
		instrmem[36] <= 32'b010001_00000_00010_0000000000000100; // m[r[0] + 4] = r[2]
		instrmem[37] <= 32'b001111_00000_00001_0000000000000011; // r[1] = m[r[0] + 3]
		instrmem[38] <= 32'b010001_00000_00001_0000000000000101; // m[r[0] + 5] = r[1]
		instrmem[39] <= 32'b001111_00000_00001_0000000000000011; // r[1] = m[r[0] + 3]
		instrmem[40] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		instrmem[41] <= 32'b010001_00000_00001_0000000000000011; // m[r[0] + 3] = r[1]
		instrmem[42] <= 32'b010100_00000000000000000000010101; // jump to 21(L2)
		instrmem[43] <= 32'b001111_00000_11101_0000000000000101; // r[29] = m[r[0] + 5]
		instrmem[44] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		instrmem[45] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[46] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[47] <= 32'b010001_00000_00001_0000000000001000; // m[r[0] + 8] = r[1]
		instrmem[48] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[49] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[50] <= 32'b010001_00000_00001_0000000000000111; // m[r[0] + 7] = r[1]
		instrmem[51] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[52] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[53] <= 32'b010001_00000_00001_0000000000000110; // m[r[0] + 6] = r[1]
		instrmem[54] <= 32'b001111_00000_00001_0000000000000111; // r[1] = m[r[0] + 7]
		instrmem[55] <= 32'b010001_00000_00001_0000000000001001; // m[r[0] + 9] = r[1]
		instrmem[56] <= 32'b001111_00000_00001_0000000000001000; // r[1] = m[r[0] + 8]
		instrmem[57] <= 32'b000011_00001_00001_0000000000000001; // r[1] = r[1] - 1
		instrmem[58] <= 32'b001111_00000_00010_0000000000001001; // r[2] = m[r[0] + 9]
		instrmem[59] <= 32'b000110_00010_00001_00101_00000_000000; // (r[2] < r[1]) ? r[5] = 1 : r[5] = 0
		instrmem[60] <= 32'b010010_00000_00101_0000000001100010; // if(r[0] == r[5]) jump to 98(L8)
		instrmem[61] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[62] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = r[a]
		instrmem[63] <= 32'b001111_00000_00001_0000000000000110; // r[1] = m[r[0] + 6]
		instrmem[64] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[65] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[66] <= 32'b001111_00000_00001_0000000000001001; // r[1] = m[r[0] + 9]
		instrmem[67] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[68] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[69] <= 32'b001111_00000_00001_0000000000001000; // r[1] = m[r[0] + 8]
		instrmem[70] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[71] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[72] <= 32'b011010_00000000000000000000000010; // jump to 2(minloc), $ra = PC + 1
		instrmem[73] <= 32'b011100_11110_11111_0000000000000000; // r[a] = stack[$sp + 0]
		instrmem[74] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[75] <= 32'b010001_00000_11101_0000000000001010; // m[r[0] + 10] = r[29]
		instrmem[76] <= 32'b001111_00000_00001_0000000000000110; // r[1] = m[r[0] + 6]
		instrmem[77] <= 32'b001111_00000_00010_0000000000001010; // r[2] = m[r[0] + 10]
		instrmem[78] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		instrmem[79] <= 32'b001111_00001_00010_0000000000000000; // r[2] = m[r[1] + 0]
		instrmem[80] <= 32'b010001_00000_00010_0000000000001011; // m[r[0] + 11] = r[2]
		instrmem[81] <= 32'b001111_00000_00001_0000000000000110; // r[1] = m[r[0] + 6]
		instrmem[82] <= 32'b001111_00000_00010_0000000000001001; // r[2] = m[r[0] + 9]
		instrmem[83] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		instrmem[84] <= 32'b001111_00000_00010_0000000000000110; // r[2] = m[r[0] + 6]
		instrmem[85] <= 32'b001111_00000_00110_0000000000001010; // r[6] = m[r[0] + 10]
		instrmem[86] <= 32'b000000_00010_00110_00010_00000_000000; // r[2] = r[2] + r[6]
		instrmem[87] <= 32'b001111_00001_00110_0000000000000000; // r[6] = m[r[1] + 0]
		instrmem[88] <= 32'b010001_00010_00110_0000000000000000; // m[r[2] + 0] = r[6]
		instrmem[89] <= 32'b001111_00000_00001_0000000000000110; // r[1] = m[r[0] + 6]
		instrmem[90] <= 32'b001111_00000_00010_0000000000001001; // r[2] = m[r[0] + 9]
		instrmem[91] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		instrmem[92] <= 32'b001111_00000_00010_0000000000001011; // r[2] = m[r[0] + 11]
		instrmem[93] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		instrmem[94] <= 32'b001111_00000_00001_0000000000001001; // r[1] = m[r[0] + 9]
		instrmem[95] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		instrmem[96] <= 32'b010001_00000_00001_0000000000001001; // m[r[0] + 9] = r[1]
		instrmem[97] <= 32'b010100_00000000000000000000111000; // jump to 56(L7)
		instrmem[98] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		instrmem[99] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[100] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[101] <= 32'b010001_00000_00001_0000000000001100; // m[r[0] + 12] = r[1]
		instrmem[102] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		instrmem[103] <= 32'b010001_00000_00001_0000000000001101; // m[r[0] + 13] = r[1]
		instrmem[104] <= 32'b001111_00000_00001_0000000000001101; // r[1] = m[r[0] + 13]
		instrmem[105] <= 32'b010000_00000_00010_0000000000000101; // r[2] = 5
		instrmem[106] <= 32'b000110_00001_00010_00110_00000_000000; // (r[1] < r[2]) ? r[6] = 1 : r[6] = 0
		instrmem[107] <= 32'b010010_00000_00110_0000000001110101; // if(r[0] == r[6]) jump to 117(L11)
		instrmem[108] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		instrmem[109] <= 32'b001111_00000_00010_0000000000001100; // r[2] = m[r[0] + 12]
		instrmem[110] <= 32'b001111_00000_00111_0000000000001101; // r[7] = m[r[0] + 13]
		instrmem[111] <= 32'b000000_00010_00111_00010_00000_000000; // r[2] = r[2] + r[7]
		instrmem[112] <= 32'b010001_00010_00001_0000000000000000; // m[r[2] + 0] = r[1]
		instrmem[113] <= 32'b001111_00000_00001_0000000000001101; // r[1] = m[r[0] + 13]
		instrmem[114] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		instrmem[115] <= 32'b010001_00000_00001_0000000000001101; // m[r[0] + 13] = r[1]
		instrmem[116] <= 32'b010100_00000000000000000001101000; // jump to 104(L10)
		instrmem[117] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		instrmem[118] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[119] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[120] <= 32'b010001_00000_00001_0000000000001111; // m[r[0] + 15] = r[1]
		instrmem[121] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[122] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[123] <= 32'b010001_00000_00001_0000000000001110; // m[r[0] + 14] = r[1]
		instrmem[124] <= 32'b001111_00000_00001_0000000000001111; // r[1] = m[r[0] + 15]
		instrmem[125] <= 32'b010000_00000_00010_0000000000000000; // r[2] = 0
		instrmem[126] <= 32'b011110_00001_00010_00111_00000_000000; // (r[1] == r[2]) ? r[7] = 1 : r[7] = 0
		instrmem[127] <= 32'b010010_00000_00111_0000000010000011; // if(r[0] == r[7]) jump to 131(L13)
		instrmem[128] <= 32'b001111_00000_11101_0000000000001110; // r[29] = m[r[0] + 14]
		instrmem[129] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		instrmem[130] <= 32'b010100_00000000000000000010010110; // jump to 150(L14)
		instrmem[131] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[132] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = r[a]
		instrmem[133] <= 32'b001111_00000_00001_0000000000001111; // r[1] = m[r[0] + 15]
		instrmem[134] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[135] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[136] <= 32'b001111_00000_00001_0000000000001110; // r[1] = m[r[0] + 14]
		instrmem[137] <= 32'b001111_00000_00010_0000000000001111; // r[2] = m[r[0] + 15]
		instrmem[138] <= 32'b001110_00001_00010_00001_00000_000000; // r[1] = r[1] / r[2]
		instrmem[139] <= 32'b001111_00000_00010_0000000000001111; // r[2] = m[r[0] + 15]
		instrmem[140] <= 32'b001101_00001_00010_00001_00000_000000; // r[1] = r[1] * r[2]
		instrmem[141] <= 32'b001111_00000_00010_0000000000001110; // r[2] = m[r[0] + 14]
		instrmem[142] <= 32'b000001_00010_00001_00010_00000_000000; // r[2] = r[2] - r[1]
		instrmem[143] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[144] <= 32'b011011_11110_00010_0000000000000000; // stack[$sp + 0] = r[2]
		instrmem[145] <= 32'b011010_00000000000000000001110110; // jump to 118(gcd), $ra = PC + 1
		instrmem[146] <= 32'b011100_11110_11111_0000000000000000; // r[a] = stack[$sp + 0]
		instrmem[147] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[148] <= 32'b000010_11101_11101_0000000000000000; // r[29] = r[29] + 0
		instrmem[149] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		instrmem[150] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[151] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[152] <= 32'b010001_00000_00001_0000000000010001; // m[r[0] + 17] = r[1]
		instrmem[153] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[154] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[155] <= 32'b010001_00000_00001_0000000000010000; // m[r[0] + 16] = r[1]
		instrmem[156] <= 32'b010000_00000_00001_0000000000000010; // r[1] = 2
		instrmem[157] <= 32'b010001_00000_00001_0000000000010010; // m[r[0] + 18] = r[1]
		instrmem[158] <= 32'b001111_00000_00001_0000000000010000; // r[1] = m[r[0] + 16]
		instrmem[159] <= 32'b000010_00001_00001_0000000000000000; // r[1] = r[1] + 0
		instrmem[160] <= 32'b010000_00000_00111_0000000000000000; // r[7] = 0
		instrmem[161] <= 32'b010001_00001_00111_0000000000000000; // m[r[1] + 0] = r[7]
		instrmem[162] <= 32'b001111_00000_00001_0000000000010000; // r[1] = m[r[0] + 16]
		instrmem[163] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		instrmem[164] <= 32'b010000_00000_00111_0000000000000001; // r[7] = 1
		instrmem[165] <= 32'b010001_00001_00111_0000000000000000; // m[r[1] + 0] = r[7]
		instrmem[166] <= 32'b001111_00000_00001_0000000000010010; // r[1] = m[r[0] + 18]
		instrmem[167] <= 32'b001111_00000_00111_0000000000010001; // r[7] = m[r[0] + 17]
		instrmem[168] <= 32'b000110_00001_00111_01000_00000_000000; // (r[1] < r[7]) ? r[8] = 1 : r[8] = 0
		instrmem[169] <= 32'b010010_00000_01000_0000000010111101; // if(r[0] == r[8]) jump to 189(L16)
		instrmem[170] <= 32'b001111_00000_00001_0000000000010010; // r[1] = m[r[0] + 18]
		instrmem[171] <= 32'b000011_00001_00001_0000000000000010; // r[1] = r[1] - 2
		instrmem[172] <= 32'b001111_00000_00111_0000000000010000; // r[7] = m[r[0] + 16]
		instrmem[173] <= 32'b000000_00111_00001_00111_00000_000000; // r[7] = r[7] + r[1]
		instrmem[174] <= 32'b001111_00000_00001_0000000000010010; // r[1] = m[r[0] + 18]
		instrmem[175] <= 32'b000011_00001_00001_0000000000000001; // r[1] = r[1] - 1
		instrmem[176] <= 32'b001111_00000_01001_0000000000010000; // r[9] = m[r[0] + 16]
		instrmem[177] <= 32'b000000_01001_00001_01001_00000_000000; // r[9] = r[9] + r[1]
		instrmem[178] <= 32'b001111_01001_00001_0000000000000000; // r[1] = m[r[9] + 0]
		instrmem[179] <= 32'b001111_00111_01010_0000000000000000; // r[10] = m[r[7] + 0]
		instrmem[180] <= 32'b000000_00001_01010_00001_00000_000000; // r[1] = r[1] + r[10]
		instrmem[181] <= 32'b001111_00000_00111_0000000000010000; // r[7] = m[r[0] + 16]
		instrmem[182] <= 32'b001111_00000_01001_0000000000010010; // r[9] = m[r[0] + 18]
		instrmem[183] <= 32'b000000_00111_01001_00111_00000_000000; // r[7] = r[7] + r[9]
		instrmem[184] <= 32'b010001_00111_00001_0000000000000000; // m[r[7] + 0] = r[1]
		instrmem[185] <= 32'b001111_00000_00001_0000000000010010; // r[1] = m[r[0] + 18]
		instrmem[186] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		instrmem[187] <= 32'b010001_00000_00001_0000000000010010; // m[r[0] + 18] = r[1]
		instrmem[188] <= 32'b010100_00000000000000000010100110; // jump to 166(L15)
		instrmem[189] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		instrmem[190] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[191] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[192] <= 32'b010001_00000_00001_0000000000010100; // m[r[0] + 20] = r[1]
		instrmem[193] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[194] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[195] <= 32'b010001_00000_00001_0000000000010011; // m[r[0] + 19] = r[1]
		instrmem[196] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		instrmem[197] <= 32'b010001_00000_00001_0000000000010101; // m[r[0] + 21] = r[1]
		instrmem[198] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		instrmem[199] <= 32'b010001_00000_00001_0000000000010110; // m[r[0] + 22] = r[1]
		instrmem[200] <= 32'b001111_00000_00001_0000000000010101; // r[1] = m[r[0] + 21]
		instrmem[201] <= 32'b001111_00000_00111_0000000000010100; // r[7] = m[r[0] + 20]
		instrmem[202] <= 32'b000110_00001_00111_01001_00000_000000; // (r[1] < r[7]) ? r[9] = 1 : r[9] = 0
		instrmem[203] <= 32'b010010_00000_01001_0000000011011100; // if(r[0] == r[9]) jump to 220(L19)
		instrmem[204] <= 32'b001111_00000_00001_0000000000010011; // r[1] = m[r[0] + 19]
		instrmem[205] <= 32'b001111_00000_00111_0000000000010101; // r[7] = m[r[0] + 21]
		instrmem[206] <= 32'b000000_00001_00111_00001_00000_000000; // r[1] = r[1] + r[7]
		instrmem[207] <= 32'b001111_00000_00111_0000000000010110; // r[7] = m[r[0] + 22]
		instrmem[208] <= 32'b001111_00001_01010_0000000000000000; // r[10] = m[r[1] + 0]
		instrmem[209] <= 32'b000110_00111_01010_00001_00000_000000; // (r[7] < r[10]) ? r[1] = 1 : r[1] = 0
		instrmem[210] <= 32'b010010_00000_00001_0000000011011000; // if(r[0] == r[1]) jump to 216(L21)
		instrmem[211] <= 32'b001111_00000_00111_0000000000010011; // r[7] = m[r[0] + 19]
		instrmem[212] <= 32'b001111_00000_01010_0000000000010101; // r[10] = m[r[0] + 21]
		instrmem[213] <= 32'b000000_00111_01010_00111_00000_000000; // r[7] = r[7] + r[10]
		instrmem[214] <= 32'b001111_00111_01010_0000000000000000; // r[10] = m[r[7] + 0]
		instrmem[215] <= 32'b010001_00000_01010_0000000000010110; // m[r[0] + 22] = r[10]
		instrmem[216] <= 32'b001111_00000_00001_0000000000010101; // r[1] = m[r[0] + 21]
		instrmem[217] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		instrmem[218] <= 32'b010001_00000_00001_0000000000010101; // m[r[0] + 21] = r[1]
		instrmem[219] <= 32'b010100_00000000000000000011001000; // jump to 200(L18)
		instrmem[220] <= 32'b001111_00000_11101_0000000000010110; // r[29] = m[r[0] + 22]
		instrmem[221] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		instrmem[222] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[223] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[224] <= 32'b010001_00000_00001_0000000000011000; // m[r[0] + 24] = r[1]
		instrmem[225] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[226] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[227] <= 32'b010001_00000_00001_0000000000010111; // m[r[0] + 23] = r[1]
		instrmem[228] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		instrmem[229] <= 32'b010001_00000_00001_0000000000011001; // m[r[0] + 25] = r[1]
		instrmem[230] <= 32'b010000_00000_00001_0000001111101000; // r[1] = 1000
		instrmem[231] <= 32'b010001_00000_00001_0000000000011010; // m[r[0] + 26] = r[1]
		instrmem[232] <= 32'b001111_00000_00001_0000000000011001; // r[1] = m[r[0] + 25]
		instrmem[233] <= 32'b001111_00000_00111_0000000000011000; // r[7] = m[r[0] + 24]
		instrmem[234] <= 32'b000110_00001_00111_01010_00000_000000; // (r[1] < r[7]) ? r[10] = 1 : r[10] = 0
		instrmem[235] <= 32'b010010_00000_01010_0000000011111100; // if(r[0] == r[10]) jump to 252(L24)
		instrmem[236] <= 32'b001111_00000_00001_0000000000010111; // r[1] = m[r[0] + 23]
		instrmem[237] <= 32'b001111_00000_00111_0000000000011001; // r[7] = m[r[0] + 25]
		instrmem[238] <= 32'b000000_00001_00111_00001_00000_000000; // r[1] = r[1] + r[7]
		instrmem[239] <= 32'b001111_00000_00111_0000000000011010; // r[7] = m[r[0] + 26]
		instrmem[240] <= 32'b001111_00001_01011_0000000000000000; // r[11] = m[r[1] + 0]
		instrmem[241] <= 32'b000110_01011_00111_00001_00000_000000; // (r[11] < r[7]) ? r[1] = 1 : r[1] = 0
		instrmem[242] <= 32'b010010_00000_00001_0000000011111000; // if(r[0] == r[1]) jump to 248(L26)
		instrmem[243] <= 32'b001111_00000_00111_0000000000010111; // r[7] = m[r[0] + 23]
		instrmem[244] <= 32'b001111_00000_01011_0000000000011001; // r[11] = m[r[0] + 25]
		instrmem[245] <= 32'b000000_00111_01011_00111_00000_000000; // r[7] = r[7] + r[11]
		instrmem[246] <= 32'b001111_00111_01011_0000000000000000; // r[11] = m[r[7] + 0]
		instrmem[247] <= 32'b010001_00000_01011_0000000000011010; // m[r[0] + 26] = r[11]
		instrmem[248] <= 32'b001111_00000_00001_0000000000011001; // r[1] = m[r[0] + 25]
		instrmem[249] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		instrmem[250] <= 32'b010001_00000_00001_0000000000011001; // m[r[0] + 25] = r[1]
		instrmem[251] <= 32'b010100_00000000000000000011101000; // jump to 232(L23)
		instrmem[252] <= 32'b001111_00000_11101_0000000000011010; // r[29] = m[r[0] + 26]
		instrmem[253] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		instrmem[254] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[255] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[256] <= 32'b010001_00000_00001_0000000000011100; // m[r[0] + 28] = r[1]
		instrmem[257] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[258] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[259] <= 32'b010001_00000_00001_0000000000011011; // m[r[0] + 27] = r[1]
		instrmem[260] <= 32'b010000_00000_00001_0000000000000001; // r[1] = 1
		instrmem[261] <= 32'b010001_00000_00001_0000000000011110; // m[r[0] + 30] = r[1]
		instrmem[262] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		instrmem[263] <= 32'b010001_00000_00001_0000000000011101; // m[r[0] + 29] = r[1]
		instrmem[264] <= 32'b001111_00000_00001_0000000000011101; // r[1] = m[r[0] + 29]
		instrmem[265] <= 32'b001111_00000_00111_0000000000011100; // r[7] = m[r[0] + 28]
		instrmem[266] <= 32'b000110_00001_00111_01011_00000_000000; // (r[1] < r[7]) ? r[11] = 1 : r[11] = 0
		instrmem[267] <= 32'b010010_00000_01011_0000000100010100; // if(r[0] == r[11]) jump to 276(L29)
		instrmem[268] <= 32'b001111_00000_00001_0000000000011110; // r[1] = m[r[0] + 30]
		instrmem[269] <= 32'b001111_00000_00111_0000000000011011; // r[7] = m[r[0] + 27]
		instrmem[270] <= 32'b001101_00001_00111_00001_00000_000000; // r[1] = r[1] * r[7]
		instrmem[271] <= 32'b010001_00000_00001_0000000000011110; // m[r[0] + 30] = r[1]
		instrmem[272] <= 32'b001111_00000_00001_0000000000011101; // r[1] = m[r[0] + 29]
		instrmem[273] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		instrmem[274] <= 32'b010001_00000_00001_0000000000011101; // m[r[0] + 29] = r[1]
		instrmem[275] <= 32'b010100_00000000000000000100001000; // jump to 264(L28)
		instrmem[276] <= 32'b001111_00000_11101_0000000000011110; // r[29] = m[r[0] + 30]
		instrmem[277] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		instrmem[278] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		instrmem[279] <= 32'b010001_00000_00001_0000000000100011; // m[r[0] + 35] = r[1]
		instrmem[280] <= 32'b001111_00000_00001_0000000000100011; // r[1] = m[r[0] + 35]
		instrmem[281] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[282] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[283] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[284] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[285] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		instrmem[286] <= 32'b001111_00000_00001_0000000000100011; // r[1] = m[r[0] + 35]
		instrmem[287] <= 32'b010000_00000_00111_0000000000000001; // r[7] = 1
		instrmem[288] <= 32'b011110_00001_00111_01100_00000_000000; // (r[1] == r[7]) ? r[12] = 1 : r[12] = 0
		instrmem[289] <= 32'b010010_00000_01100_0000000100110000; // if(r[0] == r[12]) jump to 304(L31)
		instrmem[290] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		instrmem[291] <= 32'b010001_00000_00001_0000000000100000; // m[r[0] + 32] = r[1]
		instrmem[292] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		instrmem[293] <= 32'b010001_00000_00001_0000000000100001; // m[r[0] + 33] = r[1]
		instrmem[294] <= 32'b001111_00000_00001_0000000000100001; // r[1] = m[r[0] + 33]
		instrmem[295] <= 32'b001111_00000_00111_0000000000100000; // r[7] = m[r[0] + 32]
		instrmem[296] <= 32'b000000_00001_00111_00001_00000_000000; // r[1] = r[1] + r[7]
		instrmem[297] <= 32'b010001_00000_00001_0000000000100000; // m[r[0] + 32] = r[1]
		instrmem[298] <= 32'b001111_00000_00001_0000000000100000; // r[1] = m[r[0] + 32]
		instrmem[299] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[300] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[301] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[302] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[303] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		instrmem[304] <= 32'b001111_00000_00001_0000000000100011; // r[1] = m[r[0] + 35]
		instrmem[305] <= 32'b010000_00000_00111_0000000000000010; // r[7] = 2
		instrmem[306] <= 32'b011110_00001_00111_01100_00000_000000; // (r[1] == r[7]) ? r[12] = 1 : r[12] = 0
		instrmem[307] <= 32'b010010_00000_01100_0000000101000010; // if(r[0] == r[12]) jump to 322(L33)
		instrmem[308] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		instrmem[309] <= 32'b010001_00000_00001_0000000000100000; // m[r[0] + 32] = r[1]
		instrmem[310] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		instrmem[311] <= 32'b010001_00000_00001_0000000000100001; // m[r[0] + 33] = r[1]
		instrmem[312] <= 32'b001111_00000_00001_0000000000100001; // r[1] = m[r[0] + 33]
		instrmem[313] <= 32'b001111_00000_00111_0000000000100000; // r[7] = m[r[0] + 32]
		instrmem[314] <= 32'b000001_00001_00111_00001_00000_000000; // r[1] = r[1] - r[7]
		instrmem[315] <= 32'b010001_00000_00001_0000000000100000; // m[r[0] + 32] = r[1]
		instrmem[316] <= 32'b001111_00000_00001_0000000000100000; // r[1] = m[r[0] + 32]
		instrmem[317] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[318] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[319] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[320] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[321] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		instrmem[322] <= 32'b001111_00000_00001_0000000000100011; // r[1] = m[r[0] + 35]
		instrmem[323] <= 32'b010000_00000_00111_0000000000000011; // r[7] = 3
		instrmem[324] <= 32'b011110_00001_00111_01100_00000_000000; // (r[1] == r[7]) ? r[12] = 1 : r[12] = 0
		instrmem[325] <= 32'b010010_00000_01100_0000000101010100; // if(r[0] == r[12]) jump to 340(L35)
		instrmem[326] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		instrmem[327] <= 32'b010001_00000_00001_0000000000100000; // m[r[0] + 32] = r[1]
		instrmem[328] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		instrmem[329] <= 32'b010001_00000_00001_0000000000100001; // m[r[0] + 33] = r[1]
		instrmem[330] <= 32'b001111_00000_00001_0000000000100000; // r[1] = m[r[0] + 32]
		instrmem[331] <= 32'b001111_00000_00111_0000000000100001; // r[7] = m[r[0] + 33]
		instrmem[332] <= 32'b001101_00001_00111_00001_00000_000000; // r[1] = r[1] * r[7]
		instrmem[333] <= 32'b010001_00000_00001_0000000000100000; // m[r[0] + 32] = r[1]
		instrmem[334] <= 32'b001111_00000_00001_0000000000100000; // r[1] = m[r[0] + 32]
		instrmem[335] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[336] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[337] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[338] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[339] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		instrmem[340] <= 32'b001111_00000_00001_0000000000100011; // r[1] = m[r[0] + 35]
		instrmem[341] <= 32'b010000_00000_00111_0000000000000100; // r[7] = 4
		instrmem[342] <= 32'b011110_00001_00111_01100_00000_000000; // (r[1] == r[7]) ? r[12] = 1 : r[12] = 0
		instrmem[343] <= 32'b010010_00000_01100_0000000101100110; // if(r[0] == r[12]) jump to 358(L37)
		instrmem[344] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		instrmem[345] <= 32'b010001_00000_00001_0000000000100000; // m[r[0] + 32] = r[1]
		instrmem[346] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		instrmem[347] <= 32'b010001_00000_00001_0000000000100001; // m[r[0] + 33] = r[1]
		instrmem[348] <= 32'b001111_00000_00001_0000000000100000; // r[1] = m[r[0] + 32]
		instrmem[349] <= 32'b001111_00000_00111_0000000000100001; // r[7] = m[r[0] + 33]
		instrmem[350] <= 32'b001110_00001_00111_00001_00000_000000; // r[1] = r[1] / r[7]
		instrmem[351] <= 32'b010001_00000_00001_0000000000100000; // m[r[0] + 32] = r[1]
		instrmem[352] <= 32'b001111_00000_00001_0000000000100000; // r[1] = m[r[0] + 32]
		instrmem[353] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[354] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[355] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[356] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[357] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		instrmem[358] <= 32'b001111_00000_00001_0000000000100011; // r[1] = m[r[0] + 35]
		instrmem[359] <= 32'b010000_00000_00111_0000000000000101; // r[7] = 5
		instrmem[360] <= 32'b011110_00001_00111_01100_00000_000000; // (r[1] == r[7]) ? r[12] = 1 : r[12] = 0
		instrmem[361] <= 32'b010010_00000_01100_0000000110000001; // if(r[0] == r[12]) jump to 385(L39)
		instrmem[362] <= 32'b010000_00000_00001_0000000000100101; // r[1] = 37
		instrmem[363] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[364] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[365] <= 32'b011010_00000000000000000001100011; // jump to 99(readVet), $ra = PC + 1
		instrmem[366] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		instrmem[367] <= 32'b010001_00000_00001_0000000000100100; // m[r[0] + 36] = r[1]
		instrmem[368] <= 32'b001111_00000_00001_0000000000100100; // r[1] = m[r[0] + 36]
		instrmem[369] <= 32'b010000_00000_00111_0000000000000101; // r[7] = 5
		instrmem[370] <= 32'b000110_00001_00111_01101_00000_000000; // (r[1] < r[7]) ? r[13] = 1 : r[13] = 0
		instrmem[371] <= 32'b010010_00000_01101_0000000110000001; // if(r[0] == r[13]) jump to 385(L41)
		instrmem[372] <= 32'b010000_00000_00001_0000000000100101; // r[1] = 37
		instrmem[373] <= 32'b001111_00000_00111_0000000000100100; // r[7] = m[r[0] + 36]
		instrmem[374] <= 32'b000000_00001_00111_00001_00000_000000; // r[1] = r[1] + r[7]
		instrmem[375] <= 32'b001111_00001_00111_0000000000000000; // r[7] = m[r[1] + 0]
		instrmem[376] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[377] <= 32'b011011_11110_00111_0000000000000000; // stack[$sp + 0] = r[7]
		instrmem[378] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[379] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[380] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		instrmem[381] <= 32'b001111_00000_00001_0000000000100100; // r[1] = m[r[0] + 36]
		instrmem[382] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		instrmem[383] <= 32'b010001_00000_00001_0000000000100100; // m[r[0] + 36] = r[1]
		instrmem[384] <= 32'b010100_00000000000000000101110000; // jump to 368(L40)
		instrmem[385] <= 32'b001111_00000_00001_0000000000100011; // r[1] = m[r[0] + 35]
		instrmem[386] <= 32'b010000_00000_00111_0000000000000110; // r[7] = 6
		instrmem[387] <= 32'b011110_00001_00111_01100_00000_000000; // (r[1] == r[7]) ? r[12] = 1 : r[12] = 0
		instrmem[388] <= 32'b010010_00000_01100_0000000110110100; // if(r[0] == r[12]) jump to 436(L44)
		instrmem[389] <= 32'b010000_00000_00001_0000000000100101; // r[1] = 37
		instrmem[390] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[391] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[392] <= 32'b011010_00000000000000000001100011; // jump to 99(readVet), $ra = PC + 1
		instrmem[393] <= 32'b010000_00000_00001_0000000001101111; // r[1] = 111
		instrmem[394] <= 32'b010001_00000_00001_0000000000011111; // m[r[0] + 31] = r[1]
		instrmem[395] <= 32'b010000_00000_00001_0000000000100101; // r[1] = 37
		instrmem[396] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[397] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[398] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		instrmem[399] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[400] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[401] <= 32'b010000_00000_00001_0000000000000101; // r[1] = 5
		instrmem[402] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[403] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[404] <= 32'b011010_00000000000000000000101101; // jump to 45(sort), $ra = PC + 1
		instrmem[405] <= 32'b001111_00000_00001_0000000000011111; // r[1] = m[r[0] + 31]
		instrmem[406] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[407] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[408] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[409] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[410] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		instrmem[411] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		instrmem[412] <= 32'b010001_00000_00001_0000000000100100; // m[r[0] + 36] = r[1]
		instrmem[413] <= 32'b001111_00000_00001_0000000000100100; // r[1] = m[r[0] + 36]
		instrmem[414] <= 32'b010000_00000_00111_0000000000000101; // r[7] = 5
		instrmem[415] <= 32'b000110_00001_00111_01110_00000_000000; // (r[1] < r[7]) ? r[14] = 1 : r[14] = 0
		instrmem[416] <= 32'b010010_00000_01110_0000000110101110; // if(r[0] == r[14]) jump to 430(L46)
		instrmem[417] <= 32'b010000_00000_00001_0000000000100101; // r[1] = 37
		instrmem[418] <= 32'b001111_00000_00111_0000000000100100; // r[7] = m[r[0] + 36]
		instrmem[419] <= 32'b000000_00001_00111_00001_00000_000000; // r[1] = r[1] + r[7]
		instrmem[420] <= 32'b001111_00001_00111_0000000000000000; // r[7] = m[r[1] + 0]
		instrmem[421] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[422] <= 32'b011011_11110_00111_0000000000000000; // stack[$sp + 0] = r[7]
		instrmem[423] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[424] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[425] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		instrmem[426] <= 32'b001111_00000_00001_0000000000100100; // r[1] = m[r[0] + 36]
		instrmem[427] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		instrmem[428] <= 32'b010001_00000_00001_0000000000100100; // m[r[0] + 36] = r[1]
		instrmem[429] <= 32'b010100_00000000000000000110011101; // jump to 413(L45)
		instrmem[430] <= 32'b001111_00000_00001_0000000000011111; // r[1] = m[r[0] + 31]
		instrmem[431] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[432] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[433] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[434] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[435] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		instrmem[436] <= 32'b001111_00000_00001_0000000000100011; // r[1] = m[r[0] + 35]
		instrmem[437] <= 32'b010000_00000_00111_0000000000000111; // r[7] = 7
		instrmem[438] <= 32'b011110_00001_00111_01100_00000_000000; // (r[1] == r[7]) ? r[12] = 1 : r[12] = 0
		instrmem[439] <= 32'b010010_00000_01100_0000000111001010; // if(r[0] == r[12]) jump to 458(L49)
		instrmem[440] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		instrmem[441] <= 32'b010001_00000_00001_0000000000100010; // m[r[0] + 34] = r[1]
		instrmem[442] <= 32'b010000_00000_00001_0000000000101010; // r[1] = 42
		instrmem[443] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[444] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[445] <= 32'b010000_00000_00001_0000000000001010; // r[1] = 10
		instrmem[446] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[447] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[448] <= 32'b011010_00000000000000000010010110; // jump to 150(fib), $ra = PC + 1
		instrmem[449] <= 32'b010000_00000_00001_0000000000101010; // r[1] = 42
		instrmem[450] <= 32'b001111_00000_00111_0000000000100010; // r[7] = m[r[0] + 34]
		instrmem[451] <= 32'b000000_00001_00111_00001_00000_000000; // r[1] = r[1] + r[7]
		instrmem[452] <= 32'b001111_00001_00111_0000000000000000; // r[7] = m[r[1] + 0]
		instrmem[453] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[454] <= 32'b011011_11110_00111_0000000000000000; // stack[$sp + 0] = r[7]
		instrmem[455] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[456] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[457] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		instrmem[458] <= 32'b001111_00000_00001_0000000000100011; // r[1] = m[r[0] + 35]
		instrmem[459] <= 32'b010000_00000_00111_0000000000001000; // r[7] = 8
		instrmem[460] <= 32'b011110_00001_00111_01100_00000_000000; // (r[1] == r[7]) ? r[12] = 1 : r[12] = 0
		instrmem[461] <= 32'b010010_00000_01100_0000000111100000; // if(r[0] == r[12]) jump to 480(L51)
		instrmem[462] <= 32'b010000_00000_00001_0000000000100101; // r[1] = 37
		instrmem[463] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[464] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[465] <= 32'b011010_00000000000000000001100011; // jump to 99(readVet), $ra = PC + 1
		instrmem[466] <= 32'b010000_00000_00001_0000000000100101; // r[1] = 37
		instrmem[467] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[468] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[469] <= 32'b010000_00000_00001_0000000000000101; // r[1] = 5
		instrmem[470] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[471] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[472] <= 32'b011010_00000000000000000011011110; // jump to 222(min), $ra = PC + 1
		instrmem[473] <= 32'b010001_00000_11101_0000000000100000; // m[r[0] + 32] = r[29]
		instrmem[474] <= 32'b001111_00000_00001_0000000000100000; // r[1] = m[r[0] + 32]
		instrmem[475] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[476] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[477] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[478] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[479] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		instrmem[480] <= 32'b001111_00000_00001_0000000000100011; // r[1] = m[r[0] + 35]
		instrmem[481] <= 32'b010000_00000_00111_0000000000001001; // r[7] = 9
		instrmem[482] <= 32'b011110_00001_00111_01100_00000_000000; // (r[1] == r[7]) ? r[12] = 1 : r[12] = 0
		instrmem[483] <= 32'b010010_00000_01100_0000000111110110; // if(r[0] == r[12]) jump to 502(L53)
		instrmem[484] <= 32'b010000_00000_00001_0000000000100101; // r[1] = 37
		instrmem[485] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[486] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[487] <= 32'b011010_00000000000000000001100011; // jump to 99(readVet), $ra = PC + 1
		instrmem[488] <= 32'b010000_00000_00001_0000000000100101; // r[1] = 37
		instrmem[489] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[490] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[491] <= 32'b010000_00000_00001_0000000000000101; // r[1] = 5
		instrmem[492] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[493] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[494] <= 32'b011010_00000000000000000010111110; // jump to 190(max), $ra = PC + 1
		instrmem[495] <= 32'b010001_00000_11101_0000000000100000; // m[r[0] + 32] = r[29]
		instrmem[496] <= 32'b001111_00000_00001_0000000000100000; // r[1] = m[r[0] + 32]
		instrmem[497] <= 32'b000010_11110_11110_0000000000000001; // $sp = $sp + 1
		instrmem[498] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		instrmem[499] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		instrmem[500] <= 32'b000011_11110_11110_0000000000000001; // $sp = $sp - 1
		instrmem[501] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		instrmem[502] <= 32'b010111_11111111111111111111111111; // hlt
		*/
		
