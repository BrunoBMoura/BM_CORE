/*
clk_read - auto clock
address - address for the data to be written
BIOS_out - output value for bios
*/

module BIOS
#(
	parameter DATA_WIDTH = 32, 
	parameter ADDR_WIDTH = 11
)
(
	input clk_read,
	input [(DATA_WIDTH-1):0] address,
	output reg [(DATA_WIDTH-1):0] BIOS_out
);

	reg [(DATA_WIDTH-1):0] bios_mem[(2**ADDR_WIDTH-1):0];
	initial
	begin
		bios_mem[0] <= 32'b010000_00000_11110_0000000000000000; // $sp = 0
		bios_mem[1] <= 32'b010100_00000000000000000000000010; // jump to 2(main)
		bios_mem[2] <= 32'b101000_0000000000_0000000000010110; // lcd_msg = 22
		bios_mem[3] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		bios_mem[4] <= 32'b010001_00000_00001_0000000000000011; // m[r[0] + 3] = r[1]
		bios_mem[5] <= 32'b010000_00000_00001_0000100000000000; // r[1] = 2048
		bios_mem[6] <= 32'b010001_00000_00001_0000000000000001; // m[r[0] + 1] = r[1]
		bios_mem[7] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		bios_mem[8] <= 32'b010001_00000_00001_0000000000000010; // m[r[0] + 2] = r[1]
		bios_mem[9] <= 32'b101000_0000000000_0000000000010111; // lcd_msg = 23
		bios_mem[10] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		bios_mem[11] <= 32'b010001_00000_00001_0000000000000100; // m[r[0] + 4] = r[1]
		bios_mem[12] <= 32'b001111_00000_00001_0000000000000100; // r[1] = m[r[0] + 4]
		bios_mem[13] <= 32'b010000_00000_00010_0000000000001101; // r[2] = 13
		bios_mem[14] <= 32'b011111_00001_00010_00011_00000_000000; // (r[1] != r[2]) ? r[3] = 1 : r[3] = 0
		bios_mem[15] <= 32'b010010_00000_00011_0000000000010111; // if(r[0] == r[3]) jump to 23(L3)
		bios_mem[16] <= 32'b101000_0000000000_0000000000011000; // lcd_msg = 24
		bios_mem[17] <= 32'b001111_00000_00001_0000000000000100; // r[1] = m[r[0] + 4]
		bios_mem[18] <= 32'b000010_00001_11011_0000000000000000; // r[27] = r[1] + 0
		bios_mem[19] <= 32'b101110_11011_000000000000000000000; // UART_data = LEDS = r[27]
		bios_mem[20] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		bios_mem[21] <= 32'b010001_00000_00001_0000000000000100; // m[r[0] + 4] = r[1]
		bios_mem[22] <= 32'b010100_00000000000000000000001100; // jump to 12(L2)
		bios_mem[23] <= 32'b101000_0000000000_0000000000011001; // lcd_msg = 25
		bios_mem[24] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		bios_mem[25] <= 32'b010001_00000_00001_0000000000000011; // m[r[0] + 3] = r[1]
		bios_mem[26] <= 32'b001111_00000_00001_0000000000000100; // r[1] = m[r[0] + 4]
		bios_mem[27] <= 32'b010000_00000_00010_0000000000000011; // r[2] = 3
		bios_mem[28] <= 32'b001101_00001_00010_00001_00000_000000; // r[1] = r[1] * r[2]
		bios_mem[29] <= 32'b010000_00000_00011_0000000000100111; // r[3] = 39
		bios_mem[30] <= 32'b011110_00001_00011_00100_00000_000000; // (r[1] == r[3]) ? r[4] = 1 : r[4] = 0
		bios_mem[31] <= 32'b010010_00000_00100_0000000000100011; // if(r[0] == r[4]) jump to 35(L5)
		bios_mem[32] <= 32'b101000_0000000000_0000000000011010; // lcd_msg = 26
		bios_mem[33] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		bios_mem[34] <= 32'b010001_00000_00001_0000000000000011; // m[r[0] + 3] = r[1]
		bios_mem[35] <= 32'b101000_0000000000_0000000000011011; // lcd_msg = 27
		bios_mem[36] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		bios_mem[37] <= 32'b010001_00000_00001_0000000000000011; // m[r[0] + 3] = r[1]
		bios_mem[38] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		bios_mem[39] <= 32'b010001_00000_00001_0000000000000000; // m[r[0] + 0] = r[1]
		bios_mem[40] <= 32'b001111_00000_00001_0000000000000000; // r[1] = m[r[0] + 0]
		bios_mem[41] <= 32'b001111_00000_00011_0000000000000001; // r[3] = m[r[0] + 1]
		bios_mem[42] <= 32'b000110_00001_00011_00100_00000_000000; // (r[1] < r[3]) ? r[4] = 1 : r[4] = 0
		bios_mem[43] <= 32'b010010_00000_00100_0000000000110100; // if(r[0] == r[4]) jump to 52(L8)
		bios_mem[44] <= 32'b001111_00000_00001_0000000000000010; // r[1] = m[r[0] + 2]
		bios_mem[45] <= 32'b001111_00000_00011_0000000000000000; // r[3] = m[r[0] + 0]
		bios_mem[46] <= 32'b001111_00000_00101_0000000000000000; // r[5] = m[r[0] + 0]
		bios_mem[47] <= 32'b100010_00001_00011_00101_00000000000; // mem[OS][line=r[5]] <= hd[proc=r[1]][line=r[3]]
		bios_mem[48] <= 32'b001111_00000_00001_0000000000000000; // r[1] = m[r[0] + 0]
		bios_mem[49] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		bios_mem[50] <= 32'b010001_00000_00001_0000000000000000; // m[r[0] + 0] = r[1]
		bios_mem[51] <= 32'b010100_00000000000000000000101000; // jump to 40(L7)
		bios_mem[52] <= 32'b101000_0000000000_0000000000011100; // lcd_msg = 28
		bios_mem[53] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		bios_mem[54] <= 32'b010001_00000_00001_0000000000000011; // m[r[0] + 3] = r[1]
		bios_mem[55] <= 32'b100000_00000_00000_00000_00000000000; // BIOS to Memory context
		bios_mem[56] <= 32'b010110_00000000000000000000000000; // nop
		bios_mem[57] <= 32'b111111_00000000000000000000000000; // end of the program
		bios_mem[58] <= 32'b010110_00000000000000000000000000; // nop
		bios_mem[59] <= 32'b010111_11111111111111111111111111; // hlt



	end

	always @ ( posedge clk_read )
	begin
		BIOS_out <= bios_mem[ address ];
	end

	
endmodule 




		  /*
		  bios_mem[0] <= 32'b010110_00000_00000_0000000000000000; //nop
		  bios_mem[1] <= 32'b010110_00000_00000_0000000000000000; //nop
		  bios_mem[2] <= 32'b010110_00000_00000_0000000000000000; //nop
		  bios_mem[3] <= 32'b000010_00001_00001_0000000000001010; // r[1] = r[1] + 10
		  bios_mem[4] <= 32'b000000_00001_00001_00010_00000_000000; // r[2] = r[1] + r[1]
		
		  bios_mem[5] <= 32'b101010_00000000000000000000000000; // change_read_shift
		
		  bios_mem[6] <= 32'b101001_00000000000000000000000000; //change_write_shift
		  bios_mem[7] <= 32'b000010_00001_00001_0000000000101101; // r[1] = r[1] + 45
		  bios_mem[8] <= 32'b000000_00001_00001_00010_00000_000000; // r[2] = r[1] + r[1]
		  bios_mem[9] <= 32'b101001_00000000000000000000000000; //change_write_shift
		
		  bios_mem[10] <= 32'b000000_00001_00010_00010_00000_000000; // r[2] = r[2] + r[1]
		  bios_mem[11] <= 32'b101010_00000000000000000000000000; // change_read_shift
		  bios_mem[12] <= 32'b000000_00001_00010_00011_00000_000000; // r[3] = r[1] + r[2]
		  bios_mem[13] <= 32'b000010_00011_00011_0000000000001010; // r[3] = r[3] + 10
			*/
			/*
		  bios_mem[0] <= 32'b010000_00000_11110_0000000000000000; // $sp = 0
		  bios_mem[1] <= 32'b010100_00000000000000000100010110; // jump to 278(main)
		  bios_mem[2] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[3] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[4] <= 32'b010001_00000_00001_0000000000000010; // m[r[0] + 2] = r[1]
		  bios_mem[5] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[6] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[7] <= 32'b010001_00000_00001_0000000000000001; // m[r[0] + 1] = r[1]
		  bios_mem[8] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[9] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[10] <= 32'b010001_00000_00001_0000000000000000; // m[r[0] + 0] = r[1]
		  bios_mem[11] <= 32'b001111_00000_00001_0000000000000001; // r[1] = m[r[0] + 1]
		  bios_mem[12] <= 32'b010001_00000_00001_0000000000000101; // m[r[0] + 5] = r[1]
		  bios_mem[13] <= 32'b001111_00000_00001_0000000000000000; // r[1] = m[r[0] + 0]
		  bios_mem[14] <= 32'b001111_00000_00010_0000000000000001; // r[2] = m[r[0] + 1]
		  bios_mem[15] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		  bios_mem[16] <= 32'b001111_00001_00010_0000000000000000; // r[2] = m[r[1] + 0]
		  bios_mem[17] <= 32'b010001_00000_00010_0000000000000100; // m[r[0] + 4] = r[2]
		  bios_mem[18] <= 32'b001111_00000_00001_0000000000000001; // r[1] = m[r[0] + 1]
		  bios_mem[19] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		  bios_mem[20] <= 32'b010001_00000_00001_0000000000000011; // m[r[0] + 3] = r[1]
		  bios_mem[21] <= 32'b001111_00000_00001_0000000000000011; // r[1] = m[r[0] + 3]
		  bios_mem[22] <= 32'b001111_00000_00010_0000000000000010; // r[2] = m[r[0] + 2]
		  bios_mem[23] <= 32'b000110_00001_00010_00011_00000_000000; // (r[1] < r[2]) ? r[3] = 1 : r[3] = 0
		  bios_mem[24] <= 32'b010010_00000_00011_0000000000101011; // if(r[0] == r[3]) jump to 43(L3)
		  bios_mem[25] <= 32'b001111_00000_00001_0000000000000000; // r[1] = m[r[0] + 0]
		  bios_mem[26] <= 32'b001111_00000_00010_0000000000000011; // r[2] = m[r[0] + 3]
		  bios_mem[27] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		  bios_mem[28] <= 32'b001111_00001_00010_0000000000000000; // r[2] = m[r[1] + 0]
		  bios_mem[29] <= 32'b001111_00000_00001_0000000000000100; // r[1] = m[r[0] + 4]
		  bios_mem[30] <= 32'b000110_00010_00001_00100_00000_000000; // (r[2] < r[1]) ? r[4] = 1 : r[4] = 0
		  bios_mem[31] <= 32'b010010_00000_00100_0000000000100111; // if(r[0] == r[4]) jump to 39(L5)
		  bios_mem[32] <= 32'b001111_00000_00001_0000000000000000; // r[1] = m[r[0] + 0]
		  bios_mem[33] <= 32'b001111_00000_00010_0000000000000011; // r[2] = m[r[0] + 3]
		  bios_mem[34] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		  bios_mem[35] <= 32'b001111_00001_00010_0000000000000000; // r[2] = m[r[1] + 0]
		  bios_mem[36] <= 32'b010001_00000_00010_0000000000000100; // m[r[0] + 4] = r[2]
		  bios_mem[37] <= 32'b001111_00000_00001_0000000000000011; // r[1] = m[r[0] + 3]
		  bios_mem[38] <= 32'b010001_00000_00001_0000000000000101; // m[r[0] + 5] = r[1]
		  bios_mem[39] <= 32'b001111_00000_00001_0000000000000011; // r[1] = m[r[0] + 3]
		  bios_mem[40] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		  bios_mem[41] <= 32'b010001_00000_00001_0000000000000011; // m[r[0] + 3] = r[1]
		  bios_mem[42] <= 32'b010100_00000000000000000000010101; // jump to 21(L2)
		  bios_mem[43] <= 32'b001111_00000_11101_0000000000000101; // r[29] = m[r[0] + 5]
		  bios_mem[44] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		  bios_mem[45] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[46] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[47] <= 32'b010001_00000_00001_0000000000001000; // m[r[0] + 8] = r[1]
		  bios_mem[48] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[49] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[50] <= 32'b010001_00000_00001_0000000000000111; // m[r[0] + 7] = r[1]
		  bios_mem[51] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[52] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[53] <= 32'b010001_00000_00001_0000000000000110; // m[r[0] + 6] = r[1]
		  bios_mem[54] <= 32'b001111_00000_00001_0000000000000111; // r[1] = m[r[0] + 7]
		  bios_mem[55] <= 32'b010001_00000_00001_0000000000001001; // m[r[0] + 9] = r[1]
		  bios_mem[56] <= 32'b001111_00000_00001_0000000000001000; // r[1] = m[r[0] + 8]
		  bios_mem[57] <= 32'b000011_00001_00001_0000000000000001; // r[1] = r[1] - 1
		  bios_mem[58] <= 32'b001111_00000_00010_0000000000001001; // r[2] = m[r[0] + 9]
		  bios_mem[59] <= 32'b000110_00010_00001_00100_00000_000000; // (r[2] < r[1]) ? r[4] = 1 : r[4] = 0
		  bios_mem[60] <= 32'b010010_00000_00100_0000000001100010; // if(r[0] == r[4]) jump to 98(L8)
		  bios_mem[61] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[62] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = r[a]
		  bios_mem[63] <= 32'b001111_00000_00001_0000000000000110; // r[1] = m[r[0] + 6]
		  bios_mem[64] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[65] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[66] <= 32'b001111_00000_00001_0000000000001001; // r[1] = m[r[0] + 9]
		  bios_mem[67] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[68] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[69] <= 32'b001111_00000_00001_0000000000001000; // r[1] = m[r[0] + 8]
		  bios_mem[70] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[71] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[72] <= 32'b011010_00000000000000000000000010; // jump to 2(minloc), $ra = PC + 1
		  bios_mem[73] <= 32'b011100_11110_11111_0000000000000000; // r[a] = stack[$sp + 0]
		  bios_mem[74] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[75] <= 32'b010001_00000_11101_0000000000001010; // m[r[0] + 10] = r[29]
		  bios_mem[76] <= 32'b001111_00000_00001_0000000000000110; // r[1] = m[r[0] + 6]
		  bios_mem[77] <= 32'b001111_00000_00010_0000000000001010; // r[2] = m[r[0] + 10]
		  bios_mem[78] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		  bios_mem[79] <= 32'b001111_00001_00010_0000000000000000; // r[2] = m[r[1] + 0]
		  bios_mem[80] <= 32'b010001_00000_00010_0000000000001011; // m[r[0] + 11] = r[2]
		  bios_mem[81] <= 32'b001111_00000_00001_0000000000000110; // r[1] = m[r[0] + 6]
		  bios_mem[82] <= 32'b001111_00000_00010_0000000000001001; // r[2] = m[r[0] + 9]
		  bios_mem[83] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		  bios_mem[84] <= 32'b001111_00000_00010_0000000000000110; // r[2] = m[r[0] + 6]
		  bios_mem[85] <= 32'b001111_00000_00101_0000000000001010; // r[5] = m[r[0] + 10]
		  bios_mem[86] <= 32'b000000_00010_00101_00010_00000_000000; // r[2] = r[2] + r[5]
		  bios_mem[87] <= 32'b001111_00001_00101_0000000000000000; // r[5] = m[r[1] + 0]
		  bios_mem[88] <= 32'b010001_00010_00101_0000000000000000; // m[r[2] + 0] = r[5]
		  bios_mem[89] <= 32'b001111_00000_00001_0000000000000110; // r[1] = m[r[0] + 6]
		  bios_mem[90] <= 32'b001111_00000_00010_0000000000001001; // r[2] = m[r[0] + 9]
		  bios_mem[91] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		  bios_mem[92] <= 32'b001111_00000_00010_0000000000001011; // r[2] = m[r[0] + 11]
		  bios_mem[93] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		  bios_mem[94] <= 32'b001111_00000_00001_0000000000001001; // r[1] = m[r[0] + 9]
		  bios_mem[95] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		  bios_mem[96] <= 32'b010001_00000_00001_0000000000001001; // m[r[0] + 9] = r[1]
		  bios_mem[97] <= 32'b010100_00000000000000000000111000; // jump to 56(L7)
		  bios_mem[98] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		  bios_mem[99] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[100] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[101] <= 32'b010001_00000_00001_0000000000001100; // m[r[0] + 12] = r[1]
		  bios_mem[102] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		  bios_mem[103] <= 32'b010001_00000_00001_0000000000001101; // m[r[0] + 13] = r[1]
		  bios_mem[104] <= 32'b001111_00000_00001_0000000000001101; // r[1] = m[r[0] + 13]
		  bios_mem[105] <= 32'b010000_00000_00010_0000000000000101; // r[2] = 5
		  bios_mem[106] <= 32'b000110_00001_00010_00100_00000_000000; // (r[1] < r[2]) ? r[4] = 1 : r[4] = 0
		  bios_mem[107] <= 32'b010010_00000_00100_0000000001110101; // if(r[0] == r[4]) jump to 117(L11)
		  bios_mem[108] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		  bios_mem[109] <= 32'b001111_00000_00010_0000000000001100; // r[2] = m[r[0] + 12]
		  bios_mem[110] <= 32'b001111_00000_00101_0000000000001101; // r[5] = m[r[0] + 13]
		  bios_mem[111] <= 32'b000000_00010_00101_00010_00000_000000; // r[2] = r[2] + r[5]
		  bios_mem[112] <= 32'b010001_00010_00001_0000000000000000; // m[r[2] + 0] = r[1]
		  bios_mem[113] <= 32'b001111_00000_00001_0000000000001101; // r[1] = m[r[0] + 13]
		  bios_mem[114] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		  bios_mem[115] <= 32'b010001_00000_00001_0000000000001101; // m[r[0] + 13] = r[1]
		  bios_mem[116] <= 32'b010100_00000000000000000001101000; // jump to 104(L10)
		  bios_mem[117] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		  bios_mem[118] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[119] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[120] <= 32'b010001_00000_00001_0000000000001111; // m[r[0] + 15] = r[1]
		  bios_mem[121] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[122] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[123] <= 32'b010001_00000_00001_0000000000001110; // m[r[0] + 14] = r[1]
		  bios_mem[124] <= 32'b001111_00000_00001_0000000000001111; // r[1] = m[r[0] + 15]
		  bios_mem[125] <= 32'b010000_00000_00010_0000000000000000; // r[2] = 0
		  bios_mem[126] <= 32'b011110_00001_00010_00100_00000_000000; // (r[1] == r[2]) ? r[4] = 1 : r[4] = 0
		  bios_mem[127] <= 32'b010010_00000_00100_0000000010000011; // if(r[0] == r[4]) jump to 131(L13)
		  bios_mem[128] <= 32'b001111_00000_11101_0000000000001110; // r[29] = m[r[0] + 14]
		  bios_mem[129] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		  bios_mem[130] <= 32'b010100_00000000000000000010010110; // jump to 150(L14)
		  bios_mem[131] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[132] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = r[a]
		  bios_mem[133] <= 32'b001111_00000_00001_0000000000001111; // r[1] = m[r[0] + 15]
		  bios_mem[134] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[135] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[136] <= 32'b001111_00000_00001_0000000000001110; // r[1] = m[r[0] + 14]
		  bios_mem[137] <= 32'b001111_00000_00010_0000000000001111; // r[2] = m[r[0] + 15]
		  bios_mem[138] <= 32'b001110_00001_00010_00001_00000_000000; // r[1] = r[1] / r[2]
		  bios_mem[139] <= 32'b001111_00000_00010_0000000000001111; // r[2] = m[r[0] + 15]
		  bios_mem[140] <= 32'b001101_00001_00010_00001_00000_000000; // r[1] = r[1] * r[2]
		  bios_mem[141] <= 32'b001111_00000_00010_0000000000001110; // r[2] = m[r[0] + 14]
		  bios_mem[142] <= 32'b000001_00010_00001_00010_00000_000000; // r[2] = r[2] - r[1]
		  bios_mem[143] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[144] <= 32'b011011_11110_00010_0000000000000000; // stack[$sp + 0] = r[2]
		  bios_mem[145] <= 32'b011010_00000000000000000001110110; // jump to 118(gcd), $ra = PC + 1
		  bios_mem[146] <= 32'b011100_11110_11111_0000000000000000; // r[a] = stack[$sp + 0]
		  bios_mem[147] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[148] <= 32'b000010_11101_11101_0000000000000000; // r[29] = r[29] + 0
		  bios_mem[149] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		  bios_mem[150] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[151] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[152] <= 32'b010001_00000_00001_0000000000010001; // m[r[0] + 17] = r[1]
		  bios_mem[153] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[154] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[155] <= 32'b010001_00000_00001_0000000000010000; // m[r[0] + 16] = r[1]
		  bios_mem[156] <= 32'b010000_00000_00001_0000000000000010; // r[1] = 2
		  bios_mem[157] <= 32'b010001_00000_00001_0000000000010010; // m[r[0] + 18] = r[1]
		  bios_mem[158] <= 32'b001111_00000_00001_0000000000010000; // r[1] = m[r[0] + 16]
		  bios_mem[159] <= 32'b000010_00001_00001_0000000000000000; // r[1] = r[1] + 0
		  bios_mem[160] <= 32'b010000_00000_00100_0000000000000000; // r[4] = 0
		  bios_mem[161] <= 32'b010001_00001_00100_0000000000000000; // m[r[1] + 0] = r[4]
		  bios_mem[162] <= 32'b001111_00000_00001_0000000000010000; // r[1] = m[r[0] + 16]
		  bios_mem[163] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		  bios_mem[164] <= 32'b010000_00000_00100_0000000000000001; // r[4] = 1
		  bios_mem[165] <= 32'b010001_00001_00100_0000000000000000; // m[r[1] + 0] = r[4]
		  bios_mem[166] <= 32'b001111_00000_00001_0000000000010010; // r[1] = m[r[0] + 18]
		  bios_mem[167] <= 32'b001111_00000_00100_0000000000010001; // r[4] = m[r[0] + 17]
		  bios_mem[168] <= 32'b000110_00001_00100_00101_00000_000000; // (r[1] < r[4]) ? r[5] = 1 : r[5] = 0
		  bios_mem[169] <= 32'b010010_00000_00101_0000000010111101; // if(r[0] == r[5]) jump to 189(L16)
		  bios_mem[170] <= 32'b001111_00000_00001_0000000000010010; // r[1] = m[r[0] + 18]
		  bios_mem[171] <= 32'b000011_00001_00001_0000000000000010; // r[1] = r[1] - 2
		  bios_mem[172] <= 32'b001111_00000_00100_0000000000010000; // r[4] = m[r[0] + 16]
		  bios_mem[173] <= 32'b000000_00100_00001_00100_00000_000000; // r[4] = r[4] + r[1]
		  bios_mem[174] <= 32'b001111_00000_00001_0000000000010010; // r[1] = m[r[0] + 18]
		  bios_mem[175] <= 32'b000011_00001_00001_0000000000000001; // r[1] = r[1] - 1
		  bios_mem[176] <= 32'b001111_00000_00110_0000000000010000; // r[6] = m[r[0] + 16]
		  bios_mem[177] <= 32'b000000_00110_00001_00110_00000_000000; // r[6] = r[6] + r[1]
		  bios_mem[178] <= 32'b001111_00110_00001_0000000000000000; // r[1] = m[r[6] + 0]
		  bios_mem[179] <= 32'b001111_00100_00111_0000000000000000; // r[7] = m[r[4] + 0]
		  bios_mem[180] <= 32'b000000_00001_00111_00001_00000_000000; // r[1] = r[1] + r[7]
		  bios_mem[181] <= 32'b001111_00000_00100_0000000000010000; // r[4] = m[r[0] + 16]
		  bios_mem[182] <= 32'b001111_00000_00110_0000000000010010; // r[6] = m[r[0] + 18]
		  bios_mem[183] <= 32'b000000_00100_00110_00100_00000_000000; // r[4] = r[4] + r[6]
		  bios_mem[184] <= 32'b010001_00100_00001_0000000000000000; // m[r[4] + 0] = r[1]
		  bios_mem[185] <= 32'b001111_00000_00001_0000000000010010; // r[1] = m[r[0] + 18]
		  bios_mem[186] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		  bios_mem[187] <= 32'b010001_00000_00001_0000000000010010; // m[r[0] + 18] = r[1]
		  bios_mem[188] <= 32'b010100_00000000000000000010100110; // jump to 166(L15)
		  bios_mem[189] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		  bios_mem[190] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[191] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[192] <= 32'b010001_00000_00001_0000000000010100; // m[r[0] + 20] = r[1]
		  bios_mem[193] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[194] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[195] <= 32'b010001_00000_00001_0000000000010011; // m[r[0] + 19] = r[1]
		  bios_mem[196] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		  bios_mem[197] <= 32'b010001_00000_00001_0000000000010101; // m[r[0] + 21] = r[1]
		  bios_mem[198] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		  bios_mem[199] <= 32'b010001_00000_00001_0000000000010110; // m[r[0] + 22] = r[1]
		  bios_mem[200] <= 32'b001111_00000_00001_0000000000010101; // r[1] = m[r[0] + 21]
		  bios_mem[201] <= 32'b001111_00000_00100_0000000000010100; // r[4] = m[r[0] + 20]
		  bios_mem[202] <= 32'b000110_00001_00100_00101_00000_000000; // (r[1] < r[4]) ? r[5] = 1 : r[5] = 0
		  bios_mem[203] <= 32'b010010_00000_00101_0000000011011100; // if(r[0] == r[5]) jump to 220(L19)
		  bios_mem[204] <= 32'b001111_00000_00001_0000000000010011; // r[1] = m[r[0] + 19]
		  bios_mem[205] <= 32'b001111_00000_00100_0000000000010101; // r[4] = m[r[0] + 21]
		  bios_mem[206] <= 32'b000000_00001_00100_00001_00000_000000; // r[1] = r[1] + r[4]
		  bios_mem[207] <= 32'b001111_00000_00100_0000000000010110; // r[4] = m[r[0] + 22]
		  bios_mem[208] <= 32'b001111_00001_00110_0000000000000000; // r[6] = m[r[1] + 0]
		  bios_mem[209] <= 32'b000110_00100_00110_00001_00000_000000; // (r[4] < r[6]) ? r[1] = 1 : r[1] = 0
		  bios_mem[210] <= 32'b010010_00000_00001_0000000011011000; // if(r[0] == r[1]) jump to 216(L21)
		  bios_mem[211] <= 32'b001111_00000_00100_0000000000010011; // r[4] = m[r[0] + 19]
		  bios_mem[212] <= 32'b001111_00000_00110_0000000000010101; // r[6] = m[r[0] + 21]
		  bios_mem[213] <= 32'b000000_00100_00110_00100_00000_000000; // r[4] = r[4] + r[6]
		  bios_mem[214] <= 32'b001111_00100_00110_0000000000000000; // r[6] = m[r[4] + 0]
		  bios_mem[215] <= 32'b010001_00000_00110_0000000000010110; // m[r[0] + 22] = r[6]
		  bios_mem[216] <= 32'b001111_00000_00001_0000000000010101; // r[1] = m[r[0] + 21]
		  bios_mem[217] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		  bios_mem[218] <= 32'b010001_00000_00001_0000000000010101; // m[r[0] + 21] = r[1]
		  bios_mem[219] <= 32'b010100_00000000000000000011001000; // jump to 200(L18)
		  bios_mem[220] <= 32'b001111_00000_11101_0000000000010110; // r[29] = m[r[0] + 22]
		  bios_mem[221] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		  bios_mem[222] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[223] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[224] <= 32'b010001_00000_00001_0000000000011000; // m[r[0] + 24] = r[1]
		  bios_mem[225] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[226] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[227] <= 32'b010001_00000_00001_0000000000010111; // m[r[0] + 23] = r[1]
		  bios_mem[228] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		  bios_mem[229] <= 32'b010001_00000_00001_0000000000011001; // m[r[0] + 25] = r[1]
		  bios_mem[230] <= 32'b010000_00000_00001_0000001111101000; // r[1] = 1000
		  bios_mem[231] <= 32'b010001_00000_00001_0000000000011010; // m[r[0] + 26] = r[1]
		  bios_mem[232] <= 32'b001111_00000_00001_0000000000011001; // r[1] = m[r[0] + 25]
		  bios_mem[233] <= 32'b001111_00000_00100_0000000000011000; // r[4] = m[r[0] + 24]
		  bios_mem[234] <= 32'b000110_00001_00100_00101_00000_000000; // (r[1] < r[4]) ? r[5] = 1 : r[5] = 0
		  bios_mem[235] <= 32'b010010_00000_00101_0000000011111100; // if(r[0] == r[5]) jump to 252(L24)
		  bios_mem[236] <= 32'b001111_00000_00001_0000000000010111; // r[1] = m[r[0] + 23]
		  bios_mem[237] <= 32'b001111_00000_00100_0000000000011001; // r[4] = m[r[0] + 25]
		  bios_mem[238] <= 32'b000000_00001_00100_00001_00000_000000; // r[1] = r[1] + r[4]
		  bios_mem[239] <= 32'b001111_00000_00100_0000000000011010; // r[4] = m[r[0] + 26]
		  bios_mem[240] <= 32'b001111_00001_00110_0000000000000000; // r[6] = m[r[1] + 0]
		  bios_mem[241] <= 32'b000110_00110_00100_00001_00000_000000; // (r[6] < r[4]) ? r[1] = 1 : r[1] = 0
		  bios_mem[242] <= 32'b010010_00000_00001_0000000011111000; // if(r[0] == r[1]) jump to 248(L26)
		  bios_mem[243] <= 32'b001111_00000_00100_0000000000010111; // r[4] = m[r[0] + 23]
		  bios_mem[244] <= 32'b001111_00000_00110_0000000000011001; // r[6] = m[r[0] + 25]
		  bios_mem[245] <= 32'b000000_00100_00110_00100_00000_000000; // r[4] = r[4] + r[6]
		  bios_mem[246] <= 32'b001111_00100_00110_0000000000000000; // r[6] = m[r[4] + 0]
		  bios_mem[247] <= 32'b010001_00000_00110_0000000000011010; // m[r[0] + 26] = r[6]
		  bios_mem[248] <= 32'b001111_00000_00001_0000000000011001; // r[1] = m[r[0] + 25]
		  bios_mem[249] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		  bios_mem[250] <= 32'b010001_00000_00001_0000000000011001; // m[r[0] + 25] = r[1]
		  bios_mem[251] <= 32'b010100_00000000000000000011101000; // jump to 232(L23)
		  bios_mem[252] <= 32'b001111_00000_11101_0000000000011010; // r[29] = m[r[0] + 26]
		  bios_mem[253] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		  bios_mem[254] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[255] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[256] <= 32'b010001_00000_00001_0000000000011100; // m[r[0] + 28] = r[1]
		  bios_mem[257] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[258] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[259] <= 32'b010001_00000_00001_0000000000011011; // m[r[0] + 27] = r[1]
		  bios_mem[260] <= 32'b010000_00000_00001_0000000000000001; // r[1] = 1
		  bios_mem[261] <= 32'b010001_00000_00001_0000000000011110; // m[r[0] + 30] = r[1]
		  bios_mem[262] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		  bios_mem[263] <= 32'b010001_00000_00001_0000000000011101; // m[r[0] + 29] = r[1]
		  bios_mem[264] <= 32'b001111_00000_00001_0000000000011101; // r[1] = m[r[0] + 29]
		  bios_mem[265] <= 32'b001111_00000_00100_0000000000011100; // r[4] = m[r[0] + 28]
		  bios_mem[266] <= 32'b000110_00001_00100_00101_00000_000000; // (r[1] < r[4]) ? r[5] = 1 : r[5] = 0
		  bios_mem[267] <= 32'b010010_00000_00101_0000000100010100; // if(r[0] == r[5]) jump to 276(L29)
		  bios_mem[268] <= 32'b001111_00000_00001_0000000000011110; // r[1] = m[r[0] + 30]
		  bios_mem[269] <= 32'b001111_00000_00100_0000000000011011; // r[4] = m[r[0] + 27]
		  bios_mem[270] <= 32'b001101_00001_00100_00001_00000_000000; // r[1] = r[1] * r[4]
		  bios_mem[271] <= 32'b010001_00000_00001_0000000000011110; // m[r[0] + 30] = r[1]
		  bios_mem[272] <= 32'b001111_00000_00001_0000000000011101; // r[1] = m[r[0] + 29]
		  bios_mem[273] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		  bios_mem[274] <= 32'b010001_00000_00001_0000000000011101; // m[r[0] + 29] = r[1]
		  bios_mem[275] <= 32'b010100_00000000000000000100001000; // jump to 264(L28)
		  bios_mem[276] <= 32'b001111_00000_11101_0000000000011110; // r[29] = m[r[0] + 30]
		  bios_mem[277] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		  bios_mem[278] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		  bios_mem[279] <= 32'b010001_00000_00001_0000000000100011; // m[r[0] + 35] = r[1]
		  bios_mem[280] <= 32'b001111_00000_00001_0000000000100011; // r[1] = m[r[0] + 35]
		  bios_mem[281] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[282] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[283] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[284] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[285] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		  bios_mem[286] <= 32'b001111_00000_00001_0000000000100011; // r[1] = m[r[0] + 35]
		  bios_mem[287] <= 32'b010000_00000_00100_0000000000000001; // r[4] = 1
		  bios_mem[288] <= 32'b011110_00001_00100_00101_00000_000000; // (r[1] == r[4]) ? r[5] = 1 : r[5] = 0
		  bios_mem[289] <= 32'b010010_00000_00101_0000000100110000; // if(r[0] == r[5]) jump to 304(L31)
		  bios_mem[290] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		  bios_mem[291] <= 32'b010001_00000_00001_0000000000100000; // m[r[0] + 32] = r[1]
		  bios_mem[292] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		  bios_mem[293] <= 32'b010001_00000_00001_0000000000100001; // m[r[0] + 33] = r[1]
		  bios_mem[294] <= 32'b001111_00000_00001_0000000000100001; // r[1] = m[r[0] + 33]
		  bios_mem[295] <= 32'b001111_00000_00100_0000000000100000; // r[4] = m[r[0] + 32]
		  bios_mem[296] <= 32'b000000_00001_00100_00001_00000_000000; // r[1] = r[1] + r[4]
		  bios_mem[297] <= 32'b010001_00000_00001_0000000000100000; // m[r[0] + 32] = r[1]
		  bios_mem[298] <= 32'b001111_00000_00001_0000000000100000; // r[1] = m[r[0] + 32]
		  bios_mem[299] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[300] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[301] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[302] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[303] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		  bios_mem[304] <= 32'b001111_00000_00001_0000000000100011; // r[1] = m[r[0] + 35]
		  bios_mem[305] <= 32'b010000_00000_00100_0000000000000010; // r[4] = 2
		  bios_mem[306] <= 32'b011110_00001_00100_00101_00000_000000; // (r[1] == r[4]) ? r[5] = 1 : r[5] = 0
		  bios_mem[307] <= 32'b010010_00000_00101_0000000101000010; // if(r[0] == r[5]) jump to 322(L33)
		  bios_mem[308] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		  bios_mem[309] <= 32'b010001_00000_00001_0000000000100000; // m[r[0] + 32] = r[1]
		  bios_mem[310] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		  bios_mem[311] <= 32'b010001_00000_00001_0000000000100001; // m[r[0] + 33] = r[1]
		  bios_mem[312] <= 32'b001111_00000_00001_0000000000100001; // r[1] = m[r[0] + 33]
		  bios_mem[313] <= 32'b001111_00000_00100_0000000000100000; // r[4] = m[r[0] + 32]
		  bios_mem[314] <= 32'b000001_00001_00100_00001_00000_000000; // r[1] = r[1] - r[4]
		  bios_mem[315] <= 32'b010001_00000_00001_0000000000100000; // m[r[0] + 32] = r[1]
		  bios_mem[316] <= 32'b001111_00000_00001_0000000000100000; // r[1] = m[r[0] + 32]
		  bios_mem[317] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[318] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[319] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[320] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[321] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		  bios_mem[322] <= 32'b001111_00000_00001_0000000000100011; // r[1] = m[r[0] + 35]
		  bios_mem[323] <= 32'b010000_00000_00100_0000000000000011; // r[4] = 3
		  bios_mem[324] <= 32'b011110_00001_00100_00101_00000_000000; // (r[1] == r[4]) ? r[5] = 1 : r[5] = 0
		  bios_mem[325] <= 32'b010010_00000_00101_0000000101010100; // if(r[0] == r[5]) jump to 340(L35)
		  bios_mem[326] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		  bios_mem[327] <= 32'b010001_00000_00001_0000000000100000; // m[r[0] + 32] = r[1]
		  bios_mem[328] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		  bios_mem[329] <= 32'b010001_00000_00001_0000000000100001; // m[r[0] + 33] = r[1]
		  bios_mem[330] <= 32'b001111_00000_00001_0000000000100000; // r[1] = m[r[0] + 32]
		  bios_mem[331] <= 32'b001111_00000_00100_0000000000100001; // r[4] = m[r[0] + 33]
		  bios_mem[332] <= 32'b001101_00001_00100_00001_00000_000000; // r[1] = r[1] * r[4]
		  bios_mem[333] <= 32'b010001_00000_00001_0000000000100000; // m[r[0] + 32] = r[1]
		  bios_mem[334] <= 32'b001111_00000_00001_0000000000100000; // r[1] = m[r[0] + 32]
		  bios_mem[335] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[336] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[337] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[338] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[339] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		  bios_mem[340] <= 32'b001111_00000_00001_0000000000100011; // r[1] = m[r[0] + 35]
		  bios_mem[341] <= 32'b010000_00000_00100_0000000000000100; // r[4] = 4
		  bios_mem[342] <= 32'b011110_00001_00100_00101_00000_000000; // (r[1] == r[4]) ? r[5] = 1 : r[5] = 0
		  bios_mem[343] <= 32'b010010_00000_00101_0000000101100110; // if(r[0] == r[5]) jump to 358(L37)
		  bios_mem[344] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		  bios_mem[345] <= 32'b010001_00000_00001_0000000000100000; // m[r[0] + 32] = r[1]
		  bios_mem[346] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		  bios_mem[347] <= 32'b010001_00000_00001_0000000000100001; // m[r[0] + 33] = r[1]
		  bios_mem[348] <= 32'b001111_00000_00001_0000000000100000; // r[1] = m[r[0] + 32]
		  bios_mem[349] <= 32'b001111_00000_00100_0000000000100001; // r[4] = m[r[0] + 33]
		  bios_mem[350] <= 32'b001110_00001_00100_00001_00000_000000; // r[1] = r[1] / r[4]
		  bios_mem[351] <= 32'b010001_00000_00001_0000000000100000; // m[r[0] + 32] = r[1]
		  bios_mem[352] <= 32'b001111_00000_00001_0000000000100000; // r[1] = m[r[0] + 32]
		  bios_mem[353] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[354] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[355] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[356] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[357] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		  bios_mem[358] <= 32'b001111_00000_00001_0000000000100011; // r[1] = m[r[0] + 35]
		  bios_mem[359] <= 32'b010000_00000_00100_0000000000000101; // r[4] = 5
		  bios_mem[360] <= 32'b011110_00001_00100_00101_00000_000000; // (r[1] == r[4]) ? r[5] = 1 : r[5] = 0
		  bios_mem[361] <= 32'b010010_00000_00101_0000000110000001; // if(r[0] == r[5]) jump to 385(L39)
		  bios_mem[362] <= 32'b010000_00000_00001_0000000000100101; // r[1] = 37
		  bios_mem[363] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[364] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[365] <= 32'b011010_00000000000000000001100011; // jump to 99(readVet), $ra = PC + 1
		  bios_mem[366] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		  bios_mem[367] <= 32'b010001_00000_00001_0000000000100100; // m[r[0] + 36] = r[1]
		  bios_mem[368] <= 32'b001111_00000_00001_0000000000100100; // r[1] = m[r[0] + 36]
		  bios_mem[369] <= 32'b010000_00000_00100_0000000000000101; // r[4] = 5
		  bios_mem[370] <= 32'b000110_00001_00100_00110_00000_000000; // (r[1] < r[4]) ? r[6] = 1 : r[6] = 0
		  bios_mem[371] <= 32'b010010_00000_00110_0000000110000001; // if(r[0] == r[6]) jump to 385(L41)
		  bios_mem[372] <= 32'b010000_00000_00001_0000000000100101; // r[1] = 37
		  bios_mem[373] <= 32'b001111_00000_00100_0000000000100100; // r[4] = m[r[0] + 36]
		  bios_mem[374] <= 32'b000000_00001_00100_00001_00000_000000; // r[1] = r[1] + r[4]
		  bios_mem[375] <= 32'b001111_00001_00100_0000000000000000; // r[4] = m[r[1] + 0]
		  bios_mem[376] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[377] <= 32'b011011_11110_00100_0000000000000000; // stack[$sp + 0] = r[4]
		  bios_mem[378] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[379] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[380] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		  bios_mem[381] <= 32'b001111_00000_00001_0000000000100100; // r[1] = m[r[0] + 36]
		  bios_mem[382] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		  bios_mem[383] <= 32'b010001_00000_00001_0000000000100100; // m[r[0] + 36] = r[1]
		  bios_mem[384] <= 32'b010100_00000000000000000101110000; // jump to 368(L40)
		  bios_mem[385] <= 32'b001111_00000_00001_0000000000100011; // r[1] = m[r[0] + 35]
		  bios_mem[386] <= 32'b010000_00000_00100_0000000000000110; // r[4] = 6
		  bios_mem[387] <= 32'b011110_00001_00100_00101_00000_000000; // (r[1] == r[4]) ? r[5] = 1 : r[5] = 0
		  bios_mem[388] <= 32'b010010_00000_00101_0000000110110100; // if(r[0] == r[5]) jump to 436(L44)
		  bios_mem[389] <= 32'b010000_00000_00001_0000000000100101; // r[1] = 37
		  bios_mem[390] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[391] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[392] <= 32'b011010_00000000000000000001100011; // jump to 99(readVet), $ra = PC + 1
		  bios_mem[393] <= 32'b010000_00000_00001_0000000001101111; // r[1] = 111
		  bios_mem[394] <= 32'b010001_00000_00001_0000000000011111; // m[r[0] + 31] = r[1]
		  bios_mem[395] <= 32'b010000_00000_00001_0000000000100101; // r[1] = 37
		  bios_mem[396] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[397] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[398] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		  bios_mem[399] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[400] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[401] <= 32'b010000_00000_00001_0000000000000101; // r[1] = 5
		  bios_mem[402] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[403] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[404] <= 32'b011010_00000000000000000000101101; // jump to 45(sort), $ra = PC + 1
		  bios_mem[405] <= 32'b001111_00000_00001_0000000000011111; // r[1] = m[r[0] + 31]
		  bios_mem[406] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[407] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[408] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[409] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[410] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		  bios_mem[411] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		  bios_mem[412] <= 32'b010001_00000_00001_0000000000100100; // m[r[0] + 36] = r[1]
		  bios_mem[413] <= 32'b001111_00000_00001_0000000000100100; // r[1] = m[r[0] + 36]
		  bios_mem[414] <= 32'b010000_00000_00100_0000000000000101; // r[4] = 5
		  bios_mem[415] <= 32'b000110_00001_00100_00110_00000_000000; // (r[1] < r[4]) ? r[6] = 1 : r[6] = 0
		  bios_mem[416] <= 32'b010010_00000_00110_0000000110101110; // if(r[0] == r[6]) jump to 430(L46)
		  bios_mem[417] <= 32'b010000_00000_00001_0000000000100101; // r[1] = 37
		  bios_mem[418] <= 32'b001111_00000_00100_0000000000100100; // r[4] = m[r[0] + 36]
		  bios_mem[419] <= 32'b000000_00001_00100_00001_00000_000000; // r[1] = r[1] + r[4]
		  bios_mem[420] <= 32'b001111_00001_00100_0000000000000000; // r[4] = m[r[1] + 0]
		  bios_mem[421] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[422] <= 32'b011011_11110_00100_0000000000000000; // stack[$sp + 0] = r[4]
		  bios_mem[423] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[424] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[425] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		  bios_mem[426] <= 32'b001111_00000_00001_0000000000100100; // r[1] = m[r[0] + 36]
		  bios_mem[427] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		  bios_mem[428] <= 32'b010001_00000_00001_0000000000100100; // m[r[0] + 36] = r[1]
		  bios_mem[429] <= 32'b010100_00000000000000000110011101; // jump to 413(L45)
		  bios_mem[430] <= 32'b001111_00000_00001_0000000000011111; // r[1] = m[r[0] + 31]
		  bios_mem[431] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[432] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[433] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[434] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[435] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		  bios_mem[436] <= 32'b001111_00000_00001_0000000000100011; // r[1] = m[r[0] + 35]
		  bios_mem[437] <= 32'b010000_00000_00100_0000000000000111; // r[4] = 7
		  bios_mem[438] <= 32'b011110_00001_00100_00101_00000_000000; // (r[1] == r[4]) ? r[5] = 1 : r[5] = 0
		  bios_mem[439] <= 32'b010010_00000_00101_0000000111001010; // if(r[0] == r[5]) jump to 458(L49)
		  bios_mem[440] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		  bios_mem[441] <= 32'b010001_00000_00001_0000000000100010; // m[r[0] + 34] = r[1]
		  bios_mem[442] <= 32'b010000_00000_00001_0000000000101010; // r[1] = 42
		  bios_mem[443] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[444] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[445] <= 32'b010000_00000_00001_0000000000001010; // r[1] = 10
		  bios_mem[446] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[447] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[448] <= 32'b011010_00000000000000000010010110; // jump to 150(fib), $ra = PC + 1
		  bios_mem[449] <= 32'b010000_00000_00001_0000000000101010; // r[1] = 42
		  bios_mem[450] <= 32'b001111_00000_00100_0000000000100010; // r[4] = m[r[0] + 34]
		  bios_mem[451] <= 32'b000000_00001_00100_00001_00000_000000; // r[1] = r[1] + r[4]
		  bios_mem[452] <= 32'b001111_00001_00100_0000000000000000; // r[4] = m[r[1] + 0]
		  bios_mem[453] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[454] <= 32'b011011_11110_00100_0000000000000000; // stack[$sp + 0] = r[4]
		  bios_mem[455] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[456] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[457] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		  bios_mem[458] <= 32'b001111_00000_00001_0000000000100011; // r[1] = m[r[0] + 35]
		  bios_mem[459] <= 32'b010000_00000_00100_0000000000001000; // r[4] = 8
		  bios_mem[460] <= 32'b011110_00001_00100_00101_00000_000000; // (r[1] == r[4]) ? r[5] = 1 : r[5] = 0
		  bios_mem[461] <= 32'b010010_00000_00101_0000000111100000; // if(r[0] == r[5]) jump to 480(L51)
		  bios_mem[462] <= 32'b010000_00000_00001_0000000000100101; // r[1] = 37
		  bios_mem[463] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[464] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[465] <= 32'b011010_00000000000000000001100011; // jump to 99(readVet), $ra = PC + 1
		  bios_mem[466] <= 32'b010000_00000_00001_0000000000100101; // r[1] = 37
		  bios_mem[467] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[468] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[469] <= 32'b010000_00000_00001_0000000000000101; // r[1] = 5
		  bios_mem[470] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[471] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[472] <= 32'b011010_00000000000000000011011110; // jump to 222(min), $ra = PC + 1
		  bios_mem[473] <= 32'b010001_00000_11101_0000000000100000; // m[r[0] + 32] = r[29]
		  bios_mem[474] <= 32'b001111_00000_00001_0000000000100000; // r[1] = m[r[0] + 32]
		  bios_mem[475] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[476] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[477] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[478] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[479] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		  bios_mem[480] <= 32'b001111_00000_00001_0000000000100011; // r[1] = m[r[0] + 35]
		  bios_mem[481] <= 32'b010000_00000_00100_0000000000001001; // r[4] = 9
		  bios_mem[482] <= 32'b011110_00001_00100_00101_00000_000000; // (r[1] == r[4]) ? r[5] = 1 : r[5] = 0
		  bios_mem[483] <= 32'b010010_00000_00101_0000000111110110; // if(r[0] == r[5]) jump to 502(L53)
		  bios_mem[484] <= 32'b010000_00000_00001_0000000000100101; // r[1] = 37
		  bios_mem[485] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[486] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[487] <= 32'b011010_00000000000000000001100011; // jump to 99(readVet), $ra = PC + 1
		  bios_mem[488] <= 32'b010000_00000_00001_0000000000100101; // r[1] = 37
		  bios_mem[489] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[490] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[491] <= 32'b010000_00000_00001_0000000000000101; // r[1] = 5
		  bios_mem[492] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[493] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[494] <= 32'b011010_00000000000000000010111110; // jump to 190(max), $ra = PC + 1
		  bios_mem[495] <= 32'b010001_00000_11101_0000000000100000; // m[r[0] + 32] = r[29]
		  bios_mem[496] <= 32'b001111_00000_00001_0000000000100000; // r[1] = m[r[0] + 32]
		  bios_mem[497] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		  bios_mem[498] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		  bios_mem[499] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		  bios_mem[500] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		  bios_mem[501] <= 32'b011001_00001_000000000000000000000; // LEDS = r[1]
		  bios_mem[502] <= 32'b010111_11111111111111111111111111; // hlt
		  */

/*
bios_mem[0] <= 32'b010000_00000_11110_0000000000000000; // $sp = 0
		bios_mem[1] <= 32'b010100_00000000000000000000000010; // jump to 2(main)
		bios_mem[2] <= 32'b10100000000000000000000000010110; // lcd_msg = 22
		bios_mem[3] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		bios_mem[4] <= 32'b010001_00000_00001_0000000000000011; // m[r[0] + 3] = r[1]
		bios_mem[5] <= 32'b010000_00000_00001_0000010000000000; // r[1] = 1024
		bios_mem[6] <= 32'b010001_00000_00001_0000000000000001; // m[r[0] + 1] = r[1]
		bios_mem[7] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		bios_mem[8] <= 32'b010001_00000_00001_0000000000000010; // m[r[0] + 2] = r[1]
		bios_mem[9] <= 32'b10100000000000000000000000010111; // lcd_msg = 23
		bios_mem[10] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		bios_mem[11] <= 32'b010001_00000_00001_0000000000000100; // m[r[0] + 4] = r[1]
		bios_mem[12] <= 32'b001111_00000_00001_0000000000000100; // r[1] = m[r[0] + 4]
		bios_mem[13] <= 32'b010000_00000_00010_0000000000001101; // r[2] = 13
		bios_mem[14] <= 32'b011111_00001_00010_00011_00000_000000; // (r[1] != r[2]) ? r[3] = 1 : r[3] = 0
		bios_mem[15] <= 32'b010010_00000_00011_0000000000010100; // if(r[0] == r[3]) jump to 20(L3)
		bios_mem[16] <= 32'b10100000000000000000000000011000; // lcd_msg = 24
		bios_mem[17] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		bios_mem[18] <= 32'b010001_00000_00001_0000000000000100; // m[r[0] + 4] = r[1]
		bios_mem[19] <= 32'b010100_00000000000000000000001100; // jump to 12(L2)
		bios_mem[20] <= 32'b10100000000000000000000000011001; // lcd_msg = 25
		bios_mem[21] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		bios_mem[22] <= 32'b010001_00000_00001_0000000000000011; // m[r[0] + 3] = r[1]
		bios_mem[23] <= 32'b001111_00000_00001_0000000000000100; // r[1] = m[r[0] + 4]
		bios_mem[24] <= 32'b010000_00000_00010_0000000000000011; // r[2] = 3
		bios_mem[25] <= 32'b001101_00001_00010_00001_00000_000000; // r[1] = r[1] * r[2]
		bios_mem[26] <= 32'b010000_00000_00011_0000000000100111; // r[3] = 39
		bios_mem[27] <= 32'b011110_00001_00011_00100_00000_000000; // (r[1] == r[3]) ? r[4] = 1 : r[4] = 0
		bios_mem[28] <= 32'b010010_00000_00100_0000000000100000; // if(r[0] == r[4]) jump to 32(L5)
		bios_mem[29] <= 32'b10100000000000000000000000011010; // lcd_msg = 26
		bios_mem[30] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		bios_mem[31] <= 32'b010001_00000_00001_0000000000000011; // m[r[0] + 3] = r[1]
		bios_mem[32] <= 32'b10100000000000000000000000011011; // lcd_msg = 27
		bios_mem[33] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		bios_mem[34] <= 32'b010001_00000_00001_0000000000000011; // m[r[0] + 3] = r[1]
		bios_mem[35] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		bios_mem[36] <= 32'b010001_00000_00001_0000000000000000; // m[r[0] + 0] = r[1]
		bios_mem[37] <= 32'b001111_00000_00001_0000000000000000; // r[1] = m[r[0] + 0]
		bios_mem[38] <= 32'b001111_00000_00011_0000000000000001; // r[3] = m[r[0] + 1]
		bios_mem[39] <= 32'b000110_00001_00011_00100_00000_000000; // (r[1] < r[3]) ? r[4] = 1 : r[4] = 0
		bios_mem[40] <= 32'b010010_00000_00100_0000000000110001; // if(r[0] == r[4]) jump to 49(L8)
		bios_mem[41] <= 32'b001111_00000_00001_0000000000000010; // r[1] = m[r[0] + 2]
		bios_mem[42] <= 32'b001111_00000_00011_0000000000000000; // r[3] = m[r[0] + 0]
		bios_mem[43] <= 32'b001111_00000_00101_0000000000000000; // r[5] = m[r[0] + 0]
		bios_mem[44] <= 32'b100010_00001_00011_00101_00000000000; // mem[OS][line=r[5]] <=   bios_mem[proc=r[1]][line=r[3]]
		bios_mem[45] <= 32'b001111_00000_00001_0000000000000000; // r[1] = m[r[0] + 0]
		bios_mem[46] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		bios_mem[47] <= 32'b010001_00000_00001_0000000000000000; // m[r[0] + 0] = r[1]
		bios_mem[48] <= 32'b010100_00000000000000000000100101; // jump to 37(L7)
		bios_mem[49] <= 32'b10100000000000000000000000011100; // lcd_msg = 28
		bios_mem[50] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		bios_mem[51] <= 32'b010001_00000_00001_0000000000000011; // m[r[0] + 3] = r[1]
		bios_mem[52] <= 32'b100000_00000_00000_00000_00000000000; // BIOS to Memory context
		bios_mem[53] <= 32'b010111_11111111111111111111111111; // hlt

*/
		
		
		
		
		
		
		
		
		
		/*
		  bios_mem[0] <= 32'b010110_00000_00000_0000000000000000; //nop
		  bios_mem[1] <= 32'b010110_00000_00000_0000000000000000; //nop
		  bios_mem[2] <= 32'b010110_00000_00000_0000000000000000; //nop
		  bios_mem[3] <= 32'b000010_00001_00001_0000000000001010; // r[1] = r[1] + 10
		  bios_mem[4] <= 32'b000000_00001_00001_00010_00000_000000; // r[2] = r[1] + r[1]
		
		  bios_mem[5] <= 32'b101010_00000000000000000000000000; // change_read_shift
		
		  bios_mem[6] <= 32'b101001_00000000000000000000000000; //change_write_shift
		  bios_mem[7] <= 32'b000010_00001_00001_0000000000101101; // r[1] = r[1] + 45
		  bios_mem[8] <= 32'b000000_00001_00001_00010_00000_000000; // r[2] = r[1] + r[1]
		  bios_mem[9] <= 32'b101001_00000000000000000000000000; //change_write_shift
		
		  bios_mem[10] <= 32'b000000_00001_00010_00010_00000_000000; // r[2] = r[2] + r[1]
		  bios_mem[11] <= 32'b101010_00000000000000000000000000; // change_read_shift
		  bios_mem[12] <= 32'b000000_00001_00010_00011_00000_000000; // r[3] = r[1] + r[2]
		  bios_mem[13] <= 32'b000010_00011_00011_0000000000001010; // r[3] = r[3] + 10
	*/
				
		/*
		  bios_mem[0] <= 32'b010000_00000_00011_0000000000011110; // r[3] = 30
		  bios_mem[1] <= 32'b010000_00000_00010_0000000000001111; // r[2] = 15
		  bios_mem[2] <= 32'b100111_00011_00010_00100_00000000000; // r[4] = {r[3], r[2]}
		  bios_mem[3] <= 32'b000010_00100_00100_0000000000000000; // r[4] = r[4] + 0
		*/
		/*
		  bios_mem[0] <= 32'b000010_00001_00001_0000000000000010; // r[1] = r[1] + 2
		  bios_mem[1] <= 32'b010000_00000_00011_0000000000011110; // r[3] = 30
		  bios_mem[2] <= 32'b100101_00001_00001_00011_00000000000; //   bios_mem[PROC=r[1]][line=r[1]] <= r[3]
		  bios_mem[3] <= 32'b100001_00010_000000000000000000000; // QUANTUM <= r[2]
		  bios_mem[4]	<= 32'b100100_00001_00001_00100_00000000000; // r[4] <=   bios_mem[PROC=r[1]][line=r[1]]
		  bios_mem[5] <= 32'b000010_00100_00100_0000000000001010; // r[4] = r[4] + 10
		  bios_mem[6] <= 32'b010110_00000_00000_0000000000000000; //nop
		  bios_mem[7] <= 32'b010110_00000_00000_0000000000000000; //nop
		  bios_mem[8] <= 32'b000010_00001_00001_0000000000001010; // r[1] = r[1] + 10
		*/
		/*
		  bios_mem[0] <= 32'b010000_00000_00001_0000000000001010; // r[1] = 10
		  bios_mem[1] <= 32'b100010_00000_00010_00010_00000000000; // mem[OS][line=r[2]] <=   bios_mem[proc=r[0]][line=r[2]]
		  bios_mem[2] <= 32'b000010_00010_00010_0000000000000001; // r[2] = r[2] + 1
		  bios_mem[3] <= 32'b100010_00000_00010_00010_00000000000; // mem[OS][line=r[2]] <=   bios_mem[proc=r[0]][line=r[2]]
		  bios_mem[4] <= 32'b000010_00010_00010_0000000000000001; // r[2] = r[2] + 1
		  bios_mem[5] <= 32'b100010_00000_00010_00010_00000000000; // mem[OS][line=r[2]] <=   bios_mem[proc=r[0]][line=r[2]]
		  bios_mem[6] <= 32'b000010_00010_00010_0000000000000001; // r[2] = r[2] + 1
		  bios_mem[7] <= 32'b100010_00000_00010_00010_00000000000; // mem[OS][line=r[2]] <=   bios_mem[proc=r[0]][line=r[2]]
		  bios_mem[8] <= 32'b000010_00010_00010_0000000000000001; // r[2] = r[2] + 1
		  bios_mem[9] <= 32'b100010_00000_00010_00010_00000000000; // mem[OS][line=r[2]] <=   bios_mem[proc=r[0]][line=r[2]]
		  bios_mem[10] <= 32'b000010_00010_00010_0000000000000001; // r[2] = r[2] + 1
		  bios_mem[11] <= 32'b100010_00000_00010_00010_00000000000; // mem[OS][line=r[2]] <=   bios_mem[proc=r[0]][line=r[2]]
		  bios_mem[12] <= 32'b000010_00010_00010_0000000000000001; // r[2] = r[2] + 1
		  bios_mem[13] <= 32'b100010_00000_00010_00010_00000000000; // mem[OS][line=r[2]] <=   bios_mem[proc=r[0]][line=r[2]]
		  bios_mem[14] <= 32'b100000_00000000000000000000000000; // END_BIOS
		  bios_mem[15] <= 32'b010110_00000_00000_0000000000000000; //nop
		*/
