/*
clk_read - auto clock
clk_write - divided clock
write_flag - flag used for data writing
track_line - hard drive's array index, relatively addressed with region shift
proc_num - hardware process number for region shift
input_data - data to be stored
hd_output - module output
*/

module Hard_drive
#(
	parameter DATA_WIDTH = 32, 
	parameter ADDR_WIDTH = 15, 
	parameter MAX_PROC_NUM = 16, 
	parameter REGION = (2**ADDR_WIDTH)/MAX_PROC_NUM // 2048
)
(
	input clk_read, clk_write, write_flag,
	input [(ADDR_WIDTH-1):0] track_line,
	input [(MAX_PROC_NUM-1):0] proc_num,
	input [(DATA_WIDTH-1):0] input_data, 
	output reg [(DATA_WIDTH-1):0] hd_output
);
	reg[(DATA_WIDTH-1):0] hd[(2**(ADDR_WIDTH))-1:0];
	
	initial
	begin
		//prog 0 - OS: stack = 0, mem_loc = 0
		hd[0] <= 32'b010000_00000_11110_0000000000000000; // $sp = 0
		hd[1] <= 32'b010100_00000000000000010001100110; // jump to 1126(main)
		hd[2] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[3] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[4] <= 32'b010000_00000_00001_0000000000000001; // r[1] = 1
		hd[5] <= 32'b010001_00000_00001_0000000001100001; // m[r[0] + 97] = r[1]
		hd[6] <= 32'b001111_00000_00001_0000000001100001; // r[1] = m[r[0] + 97]
		hd[7] <= 32'b001111_00000_00010_0000000000000000; // r[2] = m[r[0] + 0]
		hd[8] <= 32'b000110_00001_00010_00011_00000_000000; // (r[1] < r[2]) ? r[3] = 1 : r[3] = 0
		hd[9] <= 32'b010010_00000_00011_0000000000010011; // if(r[0] == r[3]) jump to 19(L3)
		hd[10] <= 32'b010000_00000_00001_0000000001010010; // r[1] = 82
		hd[11] <= 32'b001111_00000_00010_0000000001100001; // r[2] = m[r[0] + 97]
		hd[12] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[13] <= 32'b010000_00000_00010_0000000000000000; // r[2] = 0
		hd[14] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[15] <= 32'b001111_00000_00001_0000000001100001; // r[1] = m[r[0] + 97]
		hd[16] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[17] <= 32'b010001_00000_00001_0000000001100001; // m[r[0] + 97] = r[1]
		hd[18] <= 32'b010100_00000000000000000000000110; // jump to 6(L2)
		hd[19] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[20] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[21] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[22] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[23] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[24] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		hd[25] <= 32'b010001_00000_00001_0000000001100010; // m[r[0] + 98] = r[1]
		hd[26] <= 32'b001111_00000_00001_0000000001100010; // r[1] = m[r[0] + 98]
		hd[27] <= 32'b001111_00000_00010_0000000000000000; // r[2] = m[r[0] + 0]
		hd[28] <= 32'b000110_00001_00010_00011_00000_000000; // (r[1] < r[2]) ? r[3] = 1 : r[3] = 0
		hd[29] <= 32'b010010_00000_00011_0000000000100111; // if(r[0] == r[3]) jump to 39(L6)
		hd[30] <= 32'b010000_00000_00001_0000000001000011; // r[1] = 67
		hd[31] <= 32'b001111_00000_00010_0000000001100010; // r[2] = m[r[0] + 98]
		hd[32] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[33] <= 32'b010000_00000_00010_0000000000000000; // r[2] = 0
		hd[34] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[35] <= 32'b001111_00000_00001_0000000001100010; // r[1] = m[r[0] + 98]
		hd[36] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[37] <= 32'b010001_00000_00001_0000000001100010; // m[r[0] + 98] = r[1]
		hd[38] <= 32'b010100_00000000000000000000011010; // jump to 26(L5)
		hd[39] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[40] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[41] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[42] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[43] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[44] <= 32'b010001_00000_00001_0000000001100011; // m[r[0] + 99] = r[1]
		hd[45] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[46] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[47] <= 32'b010000_00000_00001_0000000000000001; // r[1] = 1
		hd[48] <= 32'b010001_00000_00001_0000000001100100; // m[r[0] + 100] = r[1]
		hd[49] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		hd[50] <= 32'b010001_00000_00001_0000000001100101; // m[r[0] + 101] = r[1]
		hd[51] <= 32'b001111_00000_00001_0000000001100100; // r[1] = m[r[0] + 100]
		hd[52] <= 32'b001111_00000_00010_0000000000000000; // r[2] = m[r[0] + 0]
		hd[53] <= 32'b000110_00001_00010_00011_00000_000000; // (r[1] < r[2]) ? r[3] = 1 : r[3] = 0
		hd[54] <= 32'b010010_00000_00011_0000000001000111; // if(r[0] == r[3]) jump to 71(L9)
		hd[55] <= 32'b010000_00000_00001_0000000000000111; // r[1] = 7
		hd[56] <= 32'b001111_00000_00010_0000000001100100; // r[2] = m[r[0] + 100]
		hd[57] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[58] <= 32'b001111_00001_00010_0000000000000000; // r[2] = m[r[1] + 0]
		hd[59] <= 32'b001111_00000_00001_0000000001100011; // r[1] = m[r[0] + 99]
		hd[60] <= 32'b011110_00010_00001_00100_00000_000000; // (r[2] == r[1]) ? r[4] = 1 : r[4] = 0
		hd[61] <= 32'b010010_00000_00100_0000000001000011; // if(r[0] == r[4]) jump to 67(L11)
		hd[62] <= 32'b010000_00000_00001_0000000000000001; // r[1] = 1
		hd[63] <= 32'b010001_00000_00001_0000000001100101; // m[r[0] + 101] = r[1]
		hd[64] <= 32'b001111_00000_00001_0000000000000000; // r[1] = m[r[0] + 0]
		hd[65] <= 32'b010001_00000_00001_0000000001100100; // m[r[0] + 100] = r[1]
		hd[66] <= 32'b010100_00000000000000000001000110; // jump to 70(L12)
		hd[67] <= 32'b001111_00000_00001_0000000001100100; // r[1] = m[r[0] + 100]
		hd[68] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[69] <= 32'b010001_00000_00001_0000000001100100; // m[r[0] + 100] = r[1]
		hd[70] <= 32'b010100_00000000000000000000110011; // jump to 51(L8)
		hd[71] <= 32'b001111_00000_11101_0000000001100101; // r[29] = m[r[0] + 101]
		hd[72] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[73] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[74] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[75] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[76] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[77] <= 32'b010001_00000_00001_0000000001100110; // m[r[0] + 102] = r[1]
		hd[78] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[79] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[80] <= 32'b010000_00000_00001_0000000000000001; // r[1] = 1
		hd[81] <= 32'b010001_00000_00001_0000000001100111; // m[r[0] + 103] = r[1]
		hd[82] <= 32'b001111_00000_00001_0000000001100111; // r[1] = m[r[0] + 103]
		hd[83] <= 32'b001111_00000_00010_0000000000000000; // r[2] = m[r[0] + 0]
		hd[84] <= 32'b000110_00001_00010_00011_00000_000000; // (r[1] < r[2]) ? r[3] = 1 : r[3] = 0
		hd[85] <= 32'b010010_00000_00011_0000000001100110; // if(r[0] == r[3]) jump to 102(L14)
		hd[86] <= 32'b010000_00000_00001_0000000000000111; // r[1] = 7
		hd[87] <= 32'b001111_00000_00010_0000000001100111; // r[2] = m[r[0] + 103]
		hd[88] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[89] <= 32'b001111_00001_00010_0000000000000000; // r[2] = m[r[1] + 0]
		hd[90] <= 32'b001111_00000_00001_0000000001100110; // r[1] = m[r[0] + 102]
		hd[91] <= 32'b011110_00010_00001_00100_00000_000000; // (r[2] == r[1]) ? r[4] = 1 : r[4] = 0
		hd[92] <= 32'b010010_00000_00100_0000000001100010; // if(r[0] == r[4]) jump to 98(L16)
		hd[93] <= 32'b001111_00000_00001_0000000001100111; // r[1] = m[r[0] + 103]
		hd[94] <= 32'b010001_00000_00001_0000000001101000; // m[r[0] + 104] = r[1]
		hd[95] <= 32'b001111_00000_00001_0000000000000000; // r[1] = m[r[0] + 0]
		hd[96] <= 32'b010001_00000_00001_0000000001100111; // m[r[0] + 103] = r[1]
		hd[97] <= 32'b010100_00000000000000000001100101; // jump to 101(L17)
		hd[98] <= 32'b001111_00000_00001_0000000001100111; // r[1] = m[r[0] + 103]
		hd[99] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[100] <= 32'b010001_00000_00001_0000000001100111; // m[r[0] + 103] = r[1]
		hd[101] <= 32'b010100_00000000000000000001010010; // jump to 82(L13)
		hd[102] <= 32'b001111_00000_11101_0000000001101000; // r[29] = m[r[0] + 104]
		hd[103] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[104] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[105] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[106] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[107] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[108] <= 32'b010001_00000_00001_0000000001101001; // m[r[0] + 105] = r[1]
		hd[109] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[110] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[111] <= 32'b010000_00000_00001_0000000000010110; // r[1] = 22
		hd[112] <= 32'b001111_00000_00010_0000000001101001; // r[2] = m[r[0] + 105]
		hd[113] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[114] <= 32'b010000_00000_00010_0000000000100101; // r[2] = 37
		hd[115] <= 32'b001111_00000_00011_0000000001101001; // r[3] = m[r[0] + 105]
		hd[116] <= 32'b000000_00010_00011_00010_00000_000000; // r[2] = r[2] + r[3]
		hd[117] <= 32'b001111_00010_00011_0000000000000000; // r[3] = m[r[2] + 0]
		hd[118] <= 32'b001111_00001_00100_0000000000000000; // r[4] = m[r[1] + 0]
		hd[119] <= 32'b000001_00011_00100_00011_00000_000000; // r[3] = r[3] - r[4]
		hd[120] <= 32'b010001_00000_00011_0000000001101010; // m[r[0] + 106] = r[3]
		hd[121] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		hd[122] <= 32'b010001_00000_00001_0000000001101011; // m[r[0] + 107] = r[1]
		hd[123] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[124] <= 32'b001111_00000_00010_0000000001101010; // r[2] = m[r[0] + 106]
		hd[125] <= 32'b000110_00001_00010_00011_00000_000000; // (r[1] < r[2]) ? r[3] = 1 : r[3] = 0
		hd[126] <= 32'b010010_00000_00011_0000000010000111; // if(r[0] == r[3]) jump to 135(L19)
		hd[127] <= 32'b001111_00000_00001_0000000001101001; // r[1] = m[r[0] + 105]
		hd[128] <= 32'b001111_00000_00010_0000000001101011; // r[2] = m[r[0] + 107]
		hd[129] <= 32'b001111_00000_00100_0000000001101011; // r[4] = m[r[0] + 107]
		hd[130] <= 32'b100011_00001_00010_00100_00000000000; // mem[proc=r[1]][line=r[4]] <= hd[proc=r[1]][line=r[2]]
		hd[131] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[132] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[133] <= 32'b010001_00000_00001_0000000001101011; // m[r[0] + 107] = r[1]
		hd[134] <= 32'b010100_00000000000000000001111011; // jump to 123(L18)
		hd[135] <= 32'b001111_00000_00001_0000000001101001; // r[1] = m[r[0] + 105]
		hd[136] <= 32'b001111_00000_00010_0000000000000101; // r[2] = m[r[0] + 5]
		hd[137] <= 32'b001101_00001_00010_00001_00000_000000; // r[1] = r[1] * r[2]
		hd[138] <= 32'b010001_00000_00001_0000000001101011; // m[r[0] + 107] = r[1]
		hd[139] <= 32'b001111_00000_00010_0000000001101011; // r[2] = m[r[0] + 107]
		hd[140] <= 32'b000010_00010_00010_0000000000000001; // r[2] = r[2] + 1
		hd[141] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[142] <= 32'b001111_00010_00001_0000000000000000; // r[1] = m[r[2] + 0]
		hd[143] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[144] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[145] <= 32'b000010_00001_00001_0000000000000010; // r[1] = r[1] + 2
		hd[146] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[147] <= 32'b001111_00001_00010_0000000000000000; // r[2] = m[r[1] + 0]
		hd[148] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[149] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[150] <= 32'b000010_00001_00001_0000000000000011; // r[1] = r[1] + 3
		hd[151] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[152] <= 32'b001111_00001_00011_0000000000000000; // r[3] = m[r[1] + 0]
		hd[153] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[154] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[155] <= 32'b000010_00001_00001_0000000000000100; // r[1] = r[1] + 4
		hd[156] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[157] <= 32'b001111_00001_00100_0000000000000000; // r[4] = m[r[1] + 0]
		hd[158] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[159] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[160] <= 32'b000010_00001_00001_0000000000000101; // r[1] = r[1] + 5
		hd[161] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[162] <= 32'b001111_00001_00101_0000000000000000; // r[5] = m[r[1] + 0]
		hd[163] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[164] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[165] <= 32'b000010_00001_00001_0000000000000110; // r[1] = r[1] + 6
		hd[166] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[167] <= 32'b001111_00001_00110_0000000000000000; // r[6] = m[r[1] + 0]
		hd[168] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[169] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[170] <= 32'b000010_00001_00001_0000000000000111; // r[1] = r[1] + 7
		hd[171] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[172] <= 32'b001111_00001_00111_0000000000000000; // r[7] = m[r[1] + 0]
		hd[173] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[174] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[175] <= 32'b000010_00001_00001_0000000000001000; // r[1] = r[1] + 8
		hd[176] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[177] <= 32'b001111_00001_01000_0000000000000000; // r[8] = m[r[1] + 0]
		hd[178] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[179] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[180] <= 32'b000010_00001_00001_0000000000001001; // r[1] = r[1] + 9
		hd[181] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[182] <= 32'b001111_00001_01001_0000000000000000; // r[9] = m[r[1] + 0]
		hd[183] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[184] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[185] <= 32'b000010_00001_00001_0000000000001010; // r[1] = r[1] + 10
		hd[186] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[187] <= 32'b001111_00001_01010_0000000000000000; // r[10] = m[r[1] + 0]
		hd[188] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[189] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[190] <= 32'b000010_00001_00001_0000000000001011; // r[1] = r[1] + 11
		hd[191] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[192] <= 32'b001111_00001_01011_0000000000000000; // r[11] = m[r[1] + 0]
		hd[193] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[194] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[195] <= 32'b000010_00001_00001_0000000000001100; // r[1] = r[1] + 12
		hd[196] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[197] <= 32'b001111_00001_01100_0000000000000000; // r[12] = m[r[1] + 0]
		hd[198] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[199] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[200] <= 32'b000010_00001_00001_0000000000001101; // r[1] = r[1] + 13
		hd[201] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[202] <= 32'b001111_00001_01101_0000000000000000; // r[13] = m[r[1] + 0]
		hd[203] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[204] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[205] <= 32'b000010_00001_00001_0000000000001110; // r[1] = r[1] + 14
		hd[206] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[207] <= 32'b001111_00001_01110_0000000000000000; // r[14] = m[r[1] + 0]
		hd[208] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[209] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[210] <= 32'b000010_00001_00001_0000000000001111; // r[1] = r[1] + 15
		hd[211] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[212] <= 32'b001111_00001_01111_0000000000000000; // r[15] = m[r[1] + 0]
		hd[213] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[214] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[215] <= 32'b000010_00001_00001_0000000000010000; // r[1] = r[1] + 16
		hd[216] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[217] <= 32'b001111_00001_10000_0000000000000000; // r[16] = m[r[1] + 0]
		hd[218] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[219] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[220] <= 32'b000010_00001_00001_0000000000010001; // r[1] = r[1] + 17
		hd[221] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[222] <= 32'b001111_00001_10001_0000000000000000; // r[17] = m[r[1] + 0]
		hd[223] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[224] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[225] <= 32'b000010_00001_00001_0000000000010010; // r[1] = r[1] + 18
		hd[226] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[227] <= 32'b001111_00001_10010_0000000000000000; // r[18] = m[r[1] + 0]
		hd[228] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[229] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[230] <= 32'b000010_00001_00001_0000000000010011; // r[1] = r[1] + 19
		hd[231] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[232] <= 32'b001111_00001_10011_0000000000000000; // r[19] = m[r[1] + 0]
		hd[233] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[234] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[235] <= 32'b000010_00001_00001_0000000000010100; // r[1] = r[1] + 20
		hd[236] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[237] <= 32'b001111_00001_10100_0000000000000000; // r[20] = m[r[1] + 0]
		hd[238] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[239] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[240] <= 32'b000010_00001_00001_0000000000010101; // r[1] = r[1] + 21
		hd[241] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[242] <= 32'b001111_00001_10101_0000000000000000; // r[21] = m[r[1] + 0]
		hd[243] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[244] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[245] <= 32'b000010_00001_00001_0000000000010110; // r[1] = r[1] + 22
		hd[246] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[247] <= 32'b001111_00001_10110_0000000000000000; // r[22] = m[r[1] + 0]
		hd[248] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[249] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[250] <= 32'b000010_00001_00001_0000000000010111; // r[1] = r[1] + 23
		hd[251] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[252] <= 32'b001111_00001_10111_0000000000000000; // r[23] = m[r[1] + 0]
		hd[253] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[254] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[255] <= 32'b000010_00001_00001_0000000000011000; // r[1] = r[1] + 24
		hd[256] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[257] <= 32'b001111_00001_11000_0000000000000000; // r[24] = m[r[1] + 0]
		hd[258] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[259] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[260] <= 32'b000010_00001_00001_0000000000011001; // r[1] = r[1] + 25
		hd[261] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[262] <= 32'b001111_00001_11001_0000000000000000; // r[25] = m[r[1] + 0]
		hd[263] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[264] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[265] <= 32'b000010_00001_00001_0000000000011010; // r[1] = r[1] + 26
		hd[266] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[267] <= 32'b001111_00001_11010_0000000000000000; // r[26] = m[r[1] + 0]
		hd[268] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[269] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[270] <= 32'b000010_00001_00001_0000000000011011; // r[1] = r[1] + 27
		hd[271] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[272] <= 32'b001111_00001_11011_0000000000000000; // r[27] = m[r[1] + 0]
		hd[273] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[274] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[275] <= 32'b000010_00001_00001_0000000000011100; // r[1] = r[1] + 28
		hd[276] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[277] <= 32'b001111_00001_11100_0000000000000000; // r[28] = m[r[1] + 0]
		hd[278] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[279] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[280] <= 32'b000010_00001_00001_0000000000011101; // r[1] = r[1] + 29
		hd[281] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[282] <= 32'b001111_00001_11101_0000000000000000; // r[29] = m[r[1] + 0]
		hd[283] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[284] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[285] <= 32'b000010_00001_00001_0000000000011110; // r[1] = r[1] + 30
		hd[286] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[287] <= 32'b001111_00001_11110_0000000000000000; // r[30] = m[r[1] + 0]
		hd[288] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[289] <= 32'b001111_00000_00001_0000000001101011; // r[1] = m[r[0] + 107]
		hd[290] <= 32'b000010_00001_00001_0000000000011111; // r[1] = r[1] + 31
		hd[291] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[292] <= 32'b001111_00001_11111_0000000000000000; // r[31] = m[r[1] + 0]
		hd[293] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[294] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[295] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[296] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[297] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[298] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[299] <= 32'b010001_00000_00001_0000000001101100; // m[r[0] + 108] = r[1]
		hd[300] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[301] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[302] <= 32'b001111_00000_00001_0000000001101100; // r[1] = m[r[0] + 108]
		hd[303] <= 32'b001111_00000_00010_0000000000000101; // r[2] = m[r[0] + 5]
		hd[304] <= 32'b001101_00001_00010_00001_00000_000000; // r[1] = r[1] * r[2]
		hd[305] <= 32'b010001_00000_00001_0000000001101101; // m[r[0] + 109] = r[1]
		hd[306] <= 32'b001111_00000_00010_0000000001101101; // r[2] = m[r[0] + 109]
		hd[307] <= 32'b000010_00010_00010_0000000000000001; // r[2] = r[2] + 1
		hd[308] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[309] <= 32'b000010_00001_00011_0000000000000000; // r[3] = r[1] + 0
		hd[310] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[311] <= 32'b010001_00010_00011_0000000000000000; // m[r[2] + 0] = r[3]
		hd[312] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[313] <= 32'b000010_00001_00001_0000000000000010; // r[1] = r[1] + 2
		hd[314] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[315] <= 32'b000010_00010_00011_0000000000000000; // r[3] = r[2] + 0
		hd[316] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[317] <= 32'b010001_00001_00011_0000000000000000; // m[r[1] + 0] = r[3]
		hd[318] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[319] <= 32'b000010_00001_00001_0000000000000011; // r[1] = r[1] + 3
		hd[320] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[321] <= 32'b000010_00011_00010_0000000000000000; // r[2] = r[3] + 0
		hd[322] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[323] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[324] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[325] <= 32'b000010_00001_00001_0000000000000100; // r[1] = r[1] + 4
		hd[326] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[327] <= 32'b000010_00100_00010_0000000000000000; // r[2] = r[4] + 0
		hd[328] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[329] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[330] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[331] <= 32'b000010_00001_00001_0000000000000101; // r[1] = r[1] + 5
		hd[332] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[333] <= 32'b000010_00101_00010_0000000000000000; // r[2] = r[5] + 0
		hd[334] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[335] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[336] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[337] <= 32'b000010_00001_00001_0000000000000110; // r[1] = r[1] + 6
		hd[338] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[339] <= 32'b000010_00110_00010_0000000000000000; // r[2] = r[6] + 0
		hd[340] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[341] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[342] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[343] <= 32'b000010_00001_00001_0000000000000111; // r[1] = r[1] + 7
		hd[344] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[345] <= 32'b000010_00111_00010_0000000000000000; // r[2] = r[7] + 0
		hd[346] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[347] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[348] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[349] <= 32'b000010_00001_00001_0000000000001000; // r[1] = r[1] + 8
		hd[350] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[351] <= 32'b000010_01000_00010_0000000000000000; // r[2] = r[8] + 0
		hd[352] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[353] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[354] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[355] <= 32'b000010_00001_00001_0000000000001001; // r[1] = r[1] + 9
		hd[356] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[357] <= 32'b000010_01001_00010_0000000000000000; // r[2] = r[9] + 0
		hd[358] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[359] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[360] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[361] <= 32'b000010_00001_00001_0000000000001010; // r[1] = r[1] + 10
		hd[362] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[363] <= 32'b000010_01010_00010_0000000000000000; // r[2] = r[10] + 0
		hd[364] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[365] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[366] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[367] <= 32'b000010_00001_00001_0000000000001011; // r[1] = r[1] + 11
		hd[368] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[369] <= 32'b000010_01011_00010_0000000000000000; // r[2] = r[11] + 0
		hd[370] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[371] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[372] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[373] <= 32'b000010_00001_00001_0000000000001100; // r[1] = r[1] + 12
		hd[374] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[375] <= 32'b000010_01100_00010_0000000000000000; // r[2] = r[12] + 0
		hd[376] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[377] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[378] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[379] <= 32'b000010_00001_00001_0000000000001101; // r[1] = r[1] + 13
		hd[380] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[381] <= 32'b000010_01101_00010_0000000000000000; // r[2] = r[13] + 0
		hd[382] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[383] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[384] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[385] <= 32'b000010_00001_00001_0000000000001110; // r[1] = r[1] + 14
		hd[386] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[387] <= 32'b000010_01110_00010_0000000000000000; // r[2] = r[14] + 0
		hd[388] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[389] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[390] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[391] <= 32'b000010_00001_00001_0000000000001111; // r[1] = r[1] + 15
		hd[392] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[393] <= 32'b000010_01111_00010_0000000000000000; // r[2] = r[15] + 0
		hd[394] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[395] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[396] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[397] <= 32'b000010_00001_00001_0000000000010000; // r[1] = r[1] + 16
		hd[398] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[399] <= 32'b000010_10000_00010_0000000000000000; // r[2] = r[16] + 0
		hd[400] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[401] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[402] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[403] <= 32'b000010_00001_00001_0000000000010001; // r[1] = r[1] + 17
		hd[404] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[405] <= 32'b000010_10001_00010_0000000000000000; // r[2] = r[17] + 0
		hd[406] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[407] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[408] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[409] <= 32'b000010_00001_00001_0000000000010010; // r[1] = r[1] + 18
		hd[410] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[411] <= 32'b000010_10010_00010_0000000000000000; // r[2] = r[18] + 0
		hd[412] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[413] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[414] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[415] <= 32'b000010_00001_00001_0000000000010011; // r[1] = r[1] + 19
		hd[416] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[417] <= 32'b000010_10011_00010_0000000000000000; // r[2] = r[19] + 0
		hd[418] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[419] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[420] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[421] <= 32'b000010_00001_00001_0000000000010100; // r[1] = r[1] + 20
		hd[422] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[423] <= 32'b000010_10100_00010_0000000000000000; // r[2] = r[20] + 0
		hd[424] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[425] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[426] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[427] <= 32'b000010_00001_00001_0000000000010101; // r[1] = r[1] + 21
		hd[428] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[429] <= 32'b000010_10101_00010_0000000000000000; // r[2] = r[21] + 0
		hd[430] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[431] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[432] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[433] <= 32'b000010_00001_00001_0000000000010110; // r[1] = r[1] + 22
		hd[434] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[435] <= 32'b000010_10110_00010_0000000000000000; // r[2] = r[22] + 0
		hd[436] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[437] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[438] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[439] <= 32'b000010_00001_00001_0000000000010111; // r[1] = r[1] + 23
		hd[440] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[441] <= 32'b000010_10111_00010_0000000000000000; // r[2] = r[23] + 0
		hd[442] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[443] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[444] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[445] <= 32'b000010_00001_00001_0000000000011000; // r[1] = r[1] + 24
		hd[446] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[447] <= 32'b000010_11000_00010_0000000000000000; // r[2] = r[24] + 0
		hd[448] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[449] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[450] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[451] <= 32'b000010_00001_00001_0000000000011001; // r[1] = r[1] + 25
		hd[452] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[453] <= 32'b000010_11001_00010_0000000000000000; // r[2] = r[25] + 0
		hd[454] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[455] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[456] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[457] <= 32'b000010_00001_00001_0000000000011010; // r[1] = r[1] + 26
		hd[458] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[459] <= 32'b000010_11010_00010_0000000000000000; // r[2] = r[26] + 0
		hd[460] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[461] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[462] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[463] <= 32'b000010_00001_00001_0000000000011011; // r[1] = r[1] + 27
		hd[464] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[465] <= 32'b000010_11011_00010_0000000000000000; // r[2] = r[27] + 0
		hd[466] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[467] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[468] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[469] <= 32'b000010_00001_00001_0000000000011100; // r[1] = r[1] + 28
		hd[470] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[471] <= 32'b000010_11100_00010_0000000000000000; // r[2] = r[28] + 0
		hd[472] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[473] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[474] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[475] <= 32'b000010_00001_00001_0000000000011101; // r[1] = r[1] + 29
		hd[476] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[477] <= 32'b000010_11101_00010_0000000000000000; // r[2] = r[29] + 0
		hd[478] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[479] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[480] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[481] <= 32'b000010_00001_00001_0000000000011110; // r[1] = r[1] + 30
		hd[482] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[483] <= 32'b000010_11110_00010_0000000000000000; // r[2] = r[30] + 0
		hd[484] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[485] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[486] <= 32'b001111_00000_00001_0000000001101101; // r[1] = m[r[0] + 109]
		hd[487] <= 32'b000010_00001_00001_0000000000011111; // r[1] = r[1] + 31
		hd[488] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[489] <= 32'b000010_11111_00010_0000000000000000; // r[2] = r[31] + 0
		hd[490] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[491] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[492] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[493] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[494] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[495] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[496] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[497] <= 32'b010001_00000_00001_0000000001101110; // m[r[0] + 110] = r[1]
		hd[498] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[499] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[500] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		hd[501] <= 32'b010001_00000_00001_0000000001110000; // m[r[0] + 112] = r[1]
		hd[502] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		hd[503] <= 32'b010001_00000_00001_0000000001110001; // m[r[0] + 113] = r[1]
		hd[504] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		hd[505] <= 32'b010001_00000_00001_0000000001110100; // m[r[0] + 116] = r[1]
		hd[506] <= 32'b101000_0000000000_0000000000000100; // lcd_msg = 4
		hd[507] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		hd[508] <= 32'b010001_00000_00001_0000000000000110; // m[r[0] + 6] = r[1]
		hd[509] <= 32'b001111_00000_00001_0000000001110000; // r[1] = m[r[0] + 112]
		hd[510] <= 32'b001111_00000_00010_0000000001101110; // r[2] = m[r[0] + 110]
		hd[511] <= 32'b000110_00001_00010_00011_00000_000000; // (r[1] < r[2]) ? r[3] = 1 : r[3] = 0
		hd[512] <= 32'b010010_00000_00011_0000001010000010; // if(r[0] == r[3]) jump to 642(L22)
		hd[513] <= 32'b010000_00000_00001_0000000001000011; // r[1] = 67
		hd[514] <= 32'b001111_00000_00010_0000000001110001; // r[2] = m[r[0] + 113]
		hd[515] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[516] <= 32'b001111_00001_00010_0000000000000000; // r[2] = m[r[1] + 0]
		hd[517] <= 32'b010001_00000_00010_0000000001101111; // m[r[0] + 111] = r[2]
		hd[518] <= 32'b001111_00000_00001_0000000001101111; // r[1] = m[r[0] + 111]
		hd[519] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[520] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[521] <= 32'b011010_00000000000000000001001011; // jump to 75(get_proc_idx), $ra = PC + 1
		hd[522] <= 32'b010001_00000_11101_0000000001110010; // m[r[0] + 114] = r[29]
		hd[523] <= 32'b010000_00000_00001_0000000000110100; // r[1] = 52
		hd[524] <= 32'b001111_00000_00010_0000000001110010; // r[2] = m[r[0] + 114]
		hd[525] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[526] <= 32'b001111_00001_00010_0000000000000000; // r[2] = m[r[1] + 0]
		hd[527] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		hd[528] <= 32'b011110_00010_00001_00100_00000_000000; // (r[2] == r[1]) ? r[4] = 1 : r[4] = 0
		hd[529] <= 32'b010010_00000_00100_0000001001110110; // if(r[0] == r[4]) jump to 630(L24)
		hd[530] <= 32'b010000_00000_00001_0000000001010010; // r[1] = 82
		hd[531] <= 32'b001111_00000_00010_0000000001110010; // r[2] = m[r[0] + 114]
		hd[532] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[533] <= 32'b001111_00001_00010_0000000000000000; // r[2] = m[r[1] + 0]
		hd[534] <= 32'b010001_00000_00010_0000000001110100; // m[r[0] + 116] = r[2]
		hd[535] <= 32'b001111_00000_00001_0000000001110100; // r[1] = m[r[0] + 116]
		hd[536] <= 32'b101100_00001_000000000000000000000; // process_pc = RS(r[1])
		hd[537] <= 32'b001111_00000_00001_0000000001110010; // r[1] = m[r[0] + 114]
		hd[538] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[539] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[540] <= 32'b011010_00000000000000000001101010; // jump to 106(load_proc_context), $ra = PC + 1
		hd[541] <= 32'b010110_00000000000000000000000000; // nop
		hd[542] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[543] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[544] <= 32'b001111_00000_11001_0000000001110010; // r[25] = m[r[0] + 114]
		hd[545] <= 32'b100110_11001_000000000000000000000; // process_number <= RS(r[25])
		hd[546] <= 32'b010110_00000000000000000000000000; // nop
		hd[547] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[548] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[549] <= 32'b010110_00000000000000000000000000; // nop
		hd[550] <= 32'b000010_11100_11101_0000000000000000; // r[29] = r[28] + 0
		hd[551] <= 32'b010001_00000_11101_0000000000000011; // m[r[0] + 3] = r[29]
		hd[552] <= 32'b101011_00000000000000000000000000; // r[28] = process_pc
		hd[553] <= 32'b000010_11100_11101_0000000000000000; // r[29] = r[28] + 0
		hd[554] <= 32'b010000_00000_00001_0000000001010010; // r[1] = 82
		hd[555] <= 32'b001111_00000_00010_0000000001110010; // r[2] = m[r[0] + 114]
		hd[556] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[557] <= 32'b010001_00001_11101_0000000000000000; // m[r[1] + 0] = r[29]
		hd[558] <= 32'b001111_00000_00001_0000000000000011; // r[1] = m[r[0] + 3]
		hd[559] <= 32'b010000_00000_00010_0000000000000010; // r[2] = 2
		hd[560] <= 32'b011110_00001_00010_00101_00000_000000; // (r[1] == r[2]) ? r[5] = 1 : r[5] = 0
		hd[561] <= 32'b010010_00000_00101_0000001000111100; // if(r[0] == r[5]) jump to 572(L25)
		hd[562] <= 32'b101000_0000000000_0000000000011110; // lcd_msg = 30
		hd[563] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		hd[564] <= 32'b010001_00000_00001_0000000001110011; // m[r[0] + 115] = r[1]
		hd[565] <= 32'b001111_00000_00001_0000000001110011; // r[1] = m[r[0] + 115]
		hd[566] <= 32'b000010_00001_11011_0000000000000000; // r[27] = r[1] + 0
		hd[567] <= 32'b011001_11011_000000000000000000000; // LEDS = r[27]
		hd[568] <= 32'b001111_00000_00001_0000000001110011; // r[1] = m[r[0] + 115]
		hd[569] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[570] <= 32'b000000_00001_00000_11011_00000_000000; // r[27] = r[1] + r[0]
		hd[571] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[572] <= 32'b001111_00000_00001_0000000000000011; // r[1] = m[r[0] + 3]
		hd[573] <= 32'b010000_00000_00010_0000000000000011; // r[2] = 3
		hd[574] <= 32'b011110_00001_00010_00101_00000_000000; // (r[1] == r[2]) ? r[5] = 1 : r[5] = 0
		hd[575] <= 32'b010010_00000_00101_0000001001001000; // if(r[0] == r[5]) jump to 584(L27)
		hd[576] <= 32'b101000_0000000000_0000000000011111; // lcd_msg = 31
		hd[577] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[578] <= 32'b000000_11011_00000_00001_00000_000000; // r[1] = r[27] + r[0]
		hd[579] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[580] <= 32'b010001_00000_00001_0000000001110011; // m[r[0] + 115] = r[1]
		hd[581] <= 32'b001111_00000_00001_0000000001110011; // r[1] = m[r[0] + 115]
		hd[582] <= 32'b000010_00001_11011_0000000000000000; // r[27] = r[1] + 0
		hd[583] <= 32'b011001_11011_000000000000000000000; // LEDS = r[27]
		hd[584] <= 32'b001111_00000_00001_0000000000000011; // r[1] = m[r[0] + 3]
		hd[585] <= 32'b010000_00000_00010_0000000000000100; // r[2] = 4
		hd[586] <= 32'b011110_00001_00010_00101_00000_000000; // (r[1] == r[2]) ? r[5] = 1 : r[5] = 0
		hd[587] <= 32'b010010_00000_00101_0000001001011000; // if(r[0] == r[5]) jump to 600(L29)
		hd[588] <= 32'b101000_0000000000_0000000000100000; // lcd_msg = 32
		hd[589] <= 32'b001111_00000_00001_0000000001110010; // r[1] = m[r[0] + 114]
		hd[590] <= 32'b000010_00001_11011_0000000000000000; // r[27] = r[1] + 0
		hd[591] <= 32'b011001_11011_000000000000000000000; // LEDS = r[27]
		hd[592] <= 32'b010000_00000_00001_0000000000110100; // r[1] = 52
		hd[593] <= 32'b001111_00000_00010_0000000001110010; // r[2] = m[r[0] + 114]
		hd[594] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[595] <= 32'b010000_00000_00010_0000000000000001; // r[2] = 1
		hd[596] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[597] <= 32'b001111_00000_00001_0000000001110000; // r[1] = m[r[0] + 112]
		hd[598] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[599] <= 32'b010001_00000_00001_0000000001110000; // m[r[0] + 112] = r[1]
		hd[600] <= 32'b001111_00000_00001_0000000000000011; // r[1] = m[r[0] + 3]
		hd[601] <= 32'b010000_00000_00010_0000000000000101; // r[2] = 5
		hd[602] <= 32'b011110_00001_00010_00101_00000_000000; // (r[1] == r[2]) ? r[5] = 1 : r[5] = 0
		hd[603] <= 32'b010010_00000_00101_0000001001100110; // if(r[0] == r[5]) jump to 614(L31)
		hd[604] <= 32'b101000_0000000000_0000000000100001; // lcd_msg = 33
		hd[605] <= 32'b101101_00000_00001_0000000000000000; // r[1] = UART_data
		hd[606] <= 32'b010001_00000_00001_0000000001110011; // m[r[0] + 115] = r[1]
		hd[607] <= 32'b001111_00000_00001_0000000001110011; // r[1] = m[r[0] + 115]
		hd[608] <= 32'b000010_00001_11011_0000000000000000; // r[27] = r[1] + 0
		hd[609] <= 32'b011001_11011_000000000000000000000; // LEDS = r[27]
		hd[610] <= 32'b001111_00000_00001_0000000001110011; // r[1] = m[r[0] + 115]
		hd[611] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[612] <= 32'b000000_00001_00000_11011_00000_000000; // r[27] = r[1] + r[0]
		hd[613] <= 32'b101001_00000000000000000000000000;// change registers write shift
		hd[614] <= 32'b001111_00000_00001_0000000000000011; // r[1] = m[r[0] + 3]
		hd[615] <= 32'b010000_00000_00010_0000000000000110; // r[2] = 6
		hd[616] <= 32'b011110_00001_00010_00101_00000_000000; // (r[1] == r[2]) ? r[5] = 1 : r[5] = 0
		hd[617] <= 32'b010010_00000_00101_0000001001110010; // if(r[0] == r[5]) jump to 626(L33)
		hd[618] <= 32'b101000_0000000000_0000000000100010; // lcd_msg = 34
		hd[619] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[620] <= 32'b000000_11011_00000_00001_00000_000000; // r[1] = r[27] + r[0]
		hd[621] <= 32'b101010_00000000000000000000000000; // change registers read shift
		hd[622] <= 32'b010001_00000_00001_0000000001110011; // m[r[0] + 115] = r[1]
		hd[623] <= 32'b001111_00000_00001_0000000001110011; // r[1] = m[r[0] + 115]
		hd[624] <= 32'b000010_00001_11011_0000000000000000; // r[27] = r[1] + 0
		hd[625] <= 32'b101110_11011_000000000000000000000; // UART_data = LEDS = r[27]
		hd[626] <= 32'b001111_00000_00001_0000000001110010; // r[1] = m[r[0] + 114]
		hd[627] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[628] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[629] <= 32'b011010_00000000000000000100101001; // jump to 297(store_proc_context), $ra = PC + 1
		hd[630] <= 32'b001111_00000_00001_0000000001101110; // r[1] = m[r[0] + 110]
		hd[631] <= 32'b000011_00001_00001_0000000000000001; // r[1] = r[1] - 1
		hd[632] <= 32'b001111_00000_00010_0000000001110001; // r[2] = m[r[0] + 113]
		hd[633] <= 32'b000110_00010_00001_00101_00000_000000; // (r[2] < r[1]) ? r[5] = 1 : r[5] = 0
		hd[634] <= 32'b010010_00000_00101_0000001001111111; // if(r[0] == r[5]) jump to 639(L36)
		hd[635] <= 32'b001111_00000_00001_0000000001110001; // r[1] = m[r[0] + 113]
		hd[636] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[637] <= 32'b010001_00000_00001_0000000001110001; // m[r[0] + 113] = r[1]
		hd[638] <= 32'b010100_00000000000000001010000001; // jump to 641(L37)
		hd[639] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		hd[640] <= 32'b010001_00000_00001_0000000001110001; // m[r[0] + 113] = r[1]
		hd[641] <= 32'b010100_00000000000000000111111101; // jump to 509(L21)
		hd[642] <= 32'b101000_0000000000_0000000000000101; // lcd_msg = 5
		hd[643] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		hd[644] <= 32'b010001_00000_00001_0000000000000110; // m[r[0] + 6] = r[1]
		hd[645] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[646] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[647] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[648] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[649] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[650] <= 32'b101000_0000000000_0000000000000010; // lcd_msg = 2
		hd[651] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		hd[652] <= 32'b010001_00000_00001_0000000001110101; // m[r[0] + 117] = r[1]
		hd[653] <= 32'b001111_00000_00001_0000000001110101; // r[1] = m[r[0] + 117]
		hd[654] <= 32'b000010_00001_11011_0000000000000000; // r[27] = r[1] + 0
		hd[655] <= 32'b011001_11011_000000000000000000000; // LEDS = r[27]
		hd[656] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		hd[657] <= 32'b010001_00000_00001_0000000001110110; // m[r[0] + 118] = r[1]
		hd[658] <= 32'b101000_0000000000_0000000000011101; // lcd_msg = 29
		hd[659] <= 32'b001111_00000_00001_0000000001110110; // r[1] = m[r[0] + 118]
		hd[660] <= 32'b001111_00000_00010_0000000001110101; // r[2] = m[r[0] + 117]
		hd[661] <= 32'b000110_00001_00010_00011_00000_000000; // (r[1] < r[2]) ? r[3] = 1 : r[3] = 0
		hd[662] <= 32'b010010_00000_00011_0000001010110101; // if(r[0] == r[3]) jump to 693(L39)
		hd[663] <= 32'b011000_00000_00001_0000000000000000; // r[1] = SWITCHES
		hd[664] <= 32'b010001_00000_00001_0000000001110111; // m[r[0] + 119] = r[1]
		hd[665] <= 32'b001111_00000_00001_0000000001110111; // r[1] = m[r[0] + 119]
		hd[666] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[667] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[668] <= 32'b011010_00000000000000000000101010; // jump to 42(check_ID), $ra = PC + 1
		hd[669] <= 32'b010000_00000_00010_0000000000000001; // r[2] = 1
		hd[670] <= 32'b011111_11101_00010_00101_00000_000000; // (r[29] != r[2]) ? r[5] = 1 : r[5] = 0
		hd[671] <= 32'b010010_00000_00101_0000001010100100; // if(r[0] == r[5]) jump to 676(L42)
		hd[672] <= 32'b101000_0000000000_0000000000000011; // lcd_msg = 3
		hd[673] <= 32'b011000_00000_00010_0000000000000000; // r[2] = SWITCHES
		hd[674] <= 32'b010001_00000_00010_0000000001110111; // m[r[0] + 119] = r[2]
		hd[675] <= 32'b010100_00000000000000001010011001; // jump to 665(L41)
		hd[676] <= 32'b001111_00000_00010_0000000001110111; // r[2] = m[r[0] + 119]
		hd[677] <= 32'b000010_00010_11011_0000000000000000; // r[27] = r[2] + 0
		hd[678] <= 32'b011001_11011_000000000000000000000; // LEDS = r[27]
		hd[679] <= 32'b010000_00000_00010_0000000001000011; // r[2] = 67
		hd[680] <= 32'b001111_00000_00101_0000000001110110; // r[5] = m[r[0] + 118]
		hd[681] <= 32'b000000_00010_00101_00010_00000_000000; // r[2] = r[2] + r[5]
		hd[682] <= 32'b001111_00000_00101_0000000001110111; // r[5] = m[r[0] + 119]
		hd[683] <= 32'b010001_00010_00101_0000000000000000; // m[r[2] + 0] = r[5]
		hd[684] <= 32'b010000_00000_00010_0000000000110100; // r[2] = 52
		hd[685] <= 32'b001111_00000_00101_0000000001110110; // r[5] = m[r[0] + 118]
		hd[686] <= 32'b000000_00010_00101_00010_00000_000000; // r[2] = r[2] + r[5]
		hd[687] <= 32'b010000_00000_00101_0000000000000000; // r[5] = 0
		hd[688] <= 32'b010001_00010_00101_0000000000000000; // m[r[2] + 0] = r[5]
		hd[689] <= 32'b001111_00000_00010_0000000001110110; // r[2] = m[r[0] + 118]
		hd[690] <= 32'b000010_00010_00010_0000000000000001; // r[2] = r[2] + 1
		hd[691] <= 32'b010001_00000_00010_0000000001110110; // m[r[0] + 118] = r[2]
		hd[692] <= 32'b010100_00000000000000001010010011; // jump to 659(L38)
		hd[693] <= 32'b001111_00000_00010_0000000001110101; // r[2] = m[r[0] + 117]
		hd[694] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[695] <= 32'b011011_11110_00010_0000000000000000; // stack[$sp + 0] = r[2]
		hd[696] <= 32'b011010_00000000000000000111101111; // jump to 495(round_robin), $ra = PC + 1
		hd[697] <= 32'b011010_00000000000000000000010110; // jump to 22(reset_process_queue), $ra = PC + 1
		hd[698] <= 32'b011010_00000000000000000000000010; // jump to 2(reset_program_counters), $ra = PC + 1
		hd[699] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[700] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[701] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[702] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[703] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[704] <= 32'b010000_00000_00010_0000000000000001; // r[2] = 1
		hd[705] <= 32'b010001_00000_00010_0000000001111000; // m[r[0] + 120] = r[2]
		hd[706] <= 32'b010000_00000_00010_0000000000000000; // r[2] = 0
		hd[707] <= 32'b010001_00000_00010_0000000001111001; // m[r[0] + 121] = r[2]
		hd[708] <= 32'b001111_00000_00010_0000000001111000; // r[2] = m[r[0] + 120]
		hd[709] <= 32'b001111_00000_00011_0000000000000001; // r[3] = m[r[0] + 1]
		hd[710] <= 32'b000110_00010_00011_00101_00000_000000; // (r[2] < r[3]) ? r[5] = 1 : r[5] = 0
		hd[711] <= 32'b010010_00000_00101_0000001011011000; // if(r[0] == r[5]) jump to 728(L45)
		hd[712] <= 32'b010000_00000_00010_0000000000000111; // r[2] = 7
		hd[713] <= 32'b001111_00000_00011_0000000001111000; // r[3] = m[r[0] + 120]
		hd[714] <= 32'b000000_00010_00011_00010_00000_000000; // r[2] = r[2] + r[3]
		hd[715] <= 32'b001111_00010_00011_0000000000000000; // r[3] = m[r[2] + 0]
		hd[716] <= 32'b010000_00000_00010_0000000001100011; // r[2] = 99
		hd[717] <= 32'b011110_00011_00010_00110_00000_000000; // (r[3] == r[2]) ? r[6] = 1 : r[6] = 0
		hd[718] <= 32'b010010_00000_00110_0000001011010100; // if(r[0] == r[6]) jump to 724(L47)
		hd[719] <= 32'b001111_00000_00010_0000000001111000; // r[2] = m[r[0] + 120]
		hd[720] <= 32'b010001_00000_00010_0000000001111001; // m[r[0] + 121] = r[2]
		hd[721] <= 32'b001111_00000_00010_0000000000000001; // r[2] = m[r[0] + 1]
		hd[722] <= 32'b010001_00000_00010_0000000001111000; // m[r[0] + 120] = r[2]
		hd[723] <= 32'b010100_00000000000000001011010111; // jump to 727(L48)
		hd[724] <= 32'b001111_00000_00010_0000000001111000; // r[2] = m[r[0] + 120]
		hd[725] <= 32'b000010_00010_00010_0000000000000001; // r[2] = r[2] + 1
		hd[726] <= 32'b010001_00000_00010_0000000001111000; // m[r[0] + 120] = r[2]
		hd[727] <= 32'b010100_00000000000000001011000100; // jump to 708(L44)
		hd[728] <= 32'b001111_00000_11101_0000000001111001; // r[29] = m[r[0] + 121]
		hd[729] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[730] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[731] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[732] <= 32'b011100_11110_00010_0000000000000000; // r[2] = stack[$sp + 0]
		hd[733] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[734] <= 32'b010001_00000_00010_0000000001111010; // m[r[0] + 122] = r[2]
		hd[735] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[736] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[737] <= 32'b101000_0000000000_0000000000001001; // lcd_msg = 9
		hd[738] <= 32'b011000_00000_00010_0000000000000000; // r[2] = SWITCHES
		hd[739] <= 32'b010001_00000_00010_0000000001111100; // m[r[0] + 124] = r[2]
		hd[740] <= 32'b001111_00000_00010_0000000001111100; // r[2] = m[r[0] + 124]
		hd[741] <= 32'b000010_00010_11011_0000000000000000; // r[27] = r[2] + 0
		hd[742] <= 32'b011001_11011_000000000000000000000; // LEDS = r[27]
		hd[743] <= 32'b010000_00000_00010_0000000000000000; // r[2] = 0
		hd[744] <= 32'b010001_00000_00010_0000000001111101; // m[r[0] + 125] = r[2]
		hd[745] <= 32'b001111_00000_00010_0000000001111101; // r[2] = m[r[0] + 125]
		hd[746] <= 32'b001111_00000_00011_0000000001111100; // r[3] = m[r[0] + 124]
		hd[747] <= 32'b000110_00010_00011_00101_00000_000000; // (r[2] < r[3]) ? r[5] = 1 : r[5] = 0
		hd[748] <= 32'b010010_00000_00101_0000001011111111; // if(r[0] == r[5]) jump to 767(L50)
		hd[749] <= 32'b101000_0000000000_0000000000001010; // lcd_msg = 10
		hd[750] <= 32'b011000_00000_00010_0000000000000000; // r[2] = SWITCHES
		hd[751] <= 32'b010001_00000_00010_0000000001111110; // m[r[0] + 126] = r[2]
		hd[752] <= 32'b101000_0000000000_0000000000001011; // lcd_msg = 11
		hd[753] <= 32'b011000_00000_00010_0000000000000000; // r[2] = SWITCHES
		hd[754] <= 32'b010001_00000_00010_0000000001111111; // m[r[0] + 127] = r[2]
		hd[755] <= 32'b001111_00000_00010_0000000001111110; // r[2] = m[r[0] + 126]
		hd[756] <= 32'b001111_00000_00011_0000000001111111; // r[3] = m[r[0] + 127]
		hd[757] <= 32'b100111_00010_00011_11101_00000_000000; // r[29] = {r[2],r[3]}
		hd[758] <= 32'b010001_00000_11101_0000000010000000; // m[r[0] + 128] = r[29]
		hd[759] <= 32'b001111_00000_00110_0000000001111010; // r[6] = m[r[0] + 122]
		hd[760] <= 32'b001111_00000_00111_0000000001111101; // r[7] = m[r[0] + 125]
		hd[761] <= 32'b001111_00000_01000_0000000010000000; // r[8] = m[r[0] + 128]
		hd[762] <= 32'b100101_00110_00111_01000_00000000000; // hd[proc=r[6]][line=r[7]] <= reg[8]
		hd[763] <= 32'b001111_00000_00110_0000000001111101; // r[6] = m[r[0] + 125]
		hd[764] <= 32'b000010_00110_00110_0000000000000001; // r[6] = r[6] + 1
		hd[765] <= 32'b010001_00000_00110_0000000001111101; // m[r[0] + 125] = r[6]
		hd[766] <= 32'b010100_00000000000000001011101001; // jump to 745(L49)
		hd[767] <= 32'b101000_0000000000_0000000000001100; // lcd_msg = 12
		hd[768] <= 32'b011000_00000_00101_0000000000000000; // r[5] = SWITCHES
		hd[769] <= 32'b010001_00000_00101_0000000001111011; // m[r[0] + 123] = r[5]
		hd[770] <= 32'b001111_00000_00101_0000000001111011; // r[5] = m[r[0] + 123]
		hd[771] <= 32'b000010_00101_11011_0000000000000000; // r[27] = r[5] + 0
		hd[772] <= 32'b011001_11011_000000000000000000000; // LEDS = r[27]
		hd[773] <= 32'b001111_00000_00101_0000000001111011; // r[5] = m[r[0] + 123]
		hd[774] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[775] <= 32'b011011_11110_00101_0000000000000000; // stack[$sp + 0] = r[5]
		hd[776] <= 32'b011010_00000000000000000000101010; // jump to 42(check_ID), $ra = PC + 1
		hd[777] <= 32'b010000_00000_00110_0000000000000001; // r[6] = 1
		hd[778] <= 32'b011110_11101_00110_00111_00000_000000; // (r[29] == r[6]) ? r[7] = 1 : r[7] = 0
		hd[779] <= 32'b010010_00000_00111_0000001100010000; // if(r[0] == r[7]) jump to 784(L53)
		hd[780] <= 32'b101000_0000000000_0000000000001101; // lcd_msg = 13
		hd[781] <= 32'b011000_00000_00110_0000000000000000; // r[6] = SWITCHES
		hd[782] <= 32'b010001_00000_00110_0000000001111011; // m[r[0] + 123] = r[6]
		hd[783] <= 32'b010100_00000000000000001100000101; // jump to 773(L52)
		hd[784] <= 32'b010000_00000_00110_0000000000000111; // r[6] = 7
		hd[785] <= 32'b001111_00000_00111_0000000001111010; // r[7] = m[r[0] + 122]
		hd[786] <= 32'b000000_00110_00111_00110_00000_000000; // r[6] = r[6] + r[7]
		hd[787] <= 32'b001111_00000_00111_0000000001111011; // r[7] = m[r[0] + 123]
		hd[788] <= 32'b010001_00110_00111_0000000000000000; // m[r[6] + 0] = r[7]
		hd[789] <= 32'b010000_00000_00110_0000000000010110; // r[6] = 22
		hd[790] <= 32'b001111_00000_00111_0000000001111010; // r[7] = m[r[0] + 122]
		hd[791] <= 32'b000000_00110_00111_00110_00000_000000; // r[6] = r[6] + r[7]
		hd[792] <= 32'b010000_00000_00111_0000000000000000; // r[7] = 0
		hd[793] <= 32'b010001_00110_00111_0000000000000000; // m[r[6] + 0] = r[7]
		hd[794] <= 32'b010000_00000_00110_0000000000100101; // r[6] = 37
		hd[795] <= 32'b001111_00000_00111_0000000001111010; // r[7] = m[r[0] + 122]
		hd[796] <= 32'b000000_00110_00111_00110_00000_000000; // r[6] = r[6] + r[7]
		hd[797] <= 32'b001111_00000_00111_0000000001111100; // r[7] = m[r[0] + 124]
		hd[798] <= 32'b010001_00110_00111_0000000000000000; // m[r[6] + 0] = r[7]
		hd[799] <= 32'b101000_0000000000_0000000000001110; // lcd_msg = 14
		hd[800] <= 32'b011000_00000_00110_0000000000000000; // r[6] = SWITCHES
		hd[801] <= 32'b010001_00000_00110_0000000000000110; // m[r[0] + 6] = r[6]
		hd[802] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[803] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[804] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[805] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[806] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[807] <= 32'b101000_0000000000_0000000000001111; // lcd_msg = 15
		hd[808] <= 32'b011000_00000_00110_0000000000000000; // r[6] = SWITCHES
		hd[809] <= 32'b010001_00000_00110_0000000010000010; // m[r[0] + 130] = r[6]
		hd[810] <= 32'b001111_00000_00110_0000000010000010; // r[6] = m[r[0] + 130]
		hd[811] <= 32'b000010_00110_11011_0000000000000000; // r[27] = r[6] + 0
		hd[812] <= 32'b011001_11011_000000000000000000000; // LEDS = r[27]
		hd[813] <= 32'b001111_00000_00110_0000000010000010; // r[6] = m[r[0] + 130]
		hd[814] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[815] <= 32'b011011_11110_00110_0000000000000000; // stack[$sp + 0] = r[6]
		hd[816] <= 32'b011010_00000000000000000000101010; // jump to 42(check_ID), $ra = PC + 1
		hd[817] <= 32'b010000_00000_00111_0000000000000001; // r[7] = 1
		hd[818] <= 32'b011111_11101_00111_01000_00000_000000; // (r[29] != r[7]) ? r[8] = 1 : r[8] = 0
		hd[819] <= 32'b010010_00000_01000_0000001100111000; // if(r[0] == r[8]) jump to 824(L56)
		hd[820] <= 32'b101000_0000000000_0000000000010000; // lcd_msg = 16
		hd[821] <= 32'b011000_00000_00111_0000000000000000; // r[7] = SWITCHES
		hd[822] <= 32'b010001_00000_00111_0000000010000010; // m[r[0] + 130] = r[7]
		hd[823] <= 32'b010100_00000000000000001100101101; // jump to 813(L55)
		hd[824] <= 32'b101000_0000000000_0000000000010001; // lcd_msg = 17
		hd[825] <= 32'b011000_00000_00111_0000000000000000; // r[7] = SWITCHES
		hd[826] <= 32'b010001_00000_00111_0000000010000011; // m[r[0] + 131] = r[7]
		hd[827] <= 32'b001111_00000_00111_0000000010000011; // r[7] = m[r[0] + 131]
		hd[828] <= 32'b000010_00111_11011_0000000000000000; // r[27] = r[7] + 0
		hd[829] <= 32'b011001_11011_000000000000000000000; // LEDS = r[27]
		hd[830] <= 32'b001111_00000_00111_0000000010000011; // r[7] = m[r[0] + 131]
		hd[831] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[832] <= 32'b011011_11110_00111_0000000000000000; // stack[$sp + 0] = r[7]
		hd[833] <= 32'b011010_00000000000000000000101010; // jump to 42(check_ID), $ra = PC + 1
		hd[834] <= 32'b010000_00000_01000_0000000000000001; // r[8] = 1
		hd[835] <= 32'b011110_11101_01000_01001_00000_000000; // (r[29] == r[8]) ? r[9] = 1 : r[9] = 0
		hd[836] <= 32'b010010_00000_01001_0000001101001001; // if(r[0] == r[9]) jump to 841(L59)
		hd[837] <= 32'b101000_0000000000_0000000000010010; // lcd_msg = 18
		hd[838] <= 32'b011000_00000_01000_0000000000000000; // r[8] = SWITCHES
		hd[839] <= 32'b010001_00000_01000_0000000010000011; // m[r[0] + 131] = r[8]
		hd[840] <= 32'b010100_00000000000000001100111110; // jump to 830(L58)
		hd[841] <= 32'b010000_00000_01000_0000000000000001; // r[8] = 1
		hd[842] <= 32'b010001_00000_01000_0000000010000001; // m[r[0] + 129] = r[8]
		hd[843] <= 32'b001111_00000_01000_0000000010000001; // r[8] = m[r[0] + 129]
		hd[844] <= 32'b001111_00000_01001_0000000000000000; // r[9] = m[r[0] + 0]
		hd[845] <= 32'b000110_01000_01001_01010_00000_000000; // (r[8] < r[9]) ? r[10] = 1 : r[10] = 0
		hd[846] <= 32'b010010_00000_01010_0000001101100010; // if(r[0] == r[10]) jump to 866(L62)
		hd[847] <= 32'b010000_00000_01000_0000000000000111; // r[8] = 7
		hd[848] <= 32'b001111_00000_01001_0000000010000001; // r[9] = m[r[0] + 129]
		hd[849] <= 32'b000000_01000_01001_01000_00000_000000; // r[8] = r[8] + r[9]
		hd[850] <= 32'b001111_01000_01001_0000000000000000; // r[9] = m[r[8] + 0]
		hd[851] <= 32'b001111_00000_01000_0000000010000010; // r[8] = m[r[0] + 130]
		hd[852] <= 32'b011110_01001_01000_01011_00000_000000; // (r[9] == r[8]) ? r[11] = 1 : r[11] = 0
		hd[853] <= 32'b010010_00000_01011_0000001101011110; // if(r[0] == r[11]) jump to 862(L64)
		hd[854] <= 32'b010000_00000_01000_0000000000000111; // r[8] = 7
		hd[855] <= 32'b001111_00000_01001_0000000010000001; // r[9] = m[r[0] + 129]
		hd[856] <= 32'b000000_01000_01001_01000_00000_000000; // r[8] = r[8] + r[9]
		hd[857] <= 32'b001111_00000_01001_0000000010000011; // r[9] = m[r[0] + 131]
		hd[858] <= 32'b010001_01000_01001_0000000000000000; // m[r[8] + 0] = r[9]
		hd[859] <= 32'b001111_00000_01000_0000000000000000; // r[8] = m[r[0] + 0]
		hd[860] <= 32'b010001_00000_01000_0000000010000001; // m[r[0] + 129] = r[8]
		hd[861] <= 32'b010100_00000000000000001101100001; // jump to 865(L65)
		hd[862] <= 32'b001111_00000_01000_0000000010000001; // r[8] = m[r[0] + 129]
		hd[863] <= 32'b000010_01000_01000_0000000000000001; // r[8] = r[8] + 1
		hd[864] <= 32'b010001_00000_01000_0000000010000001; // m[r[0] + 129] = r[8]
		hd[865] <= 32'b010100_00000000000000001101001011; // jump to 843(L61)
		hd[866] <= 32'b101000_0000000000_0000000000010011; // lcd_msg = 19
		hd[867] <= 32'b011000_00000_01000_0000000000000000; // r[8] = SWITCHES
		hd[868] <= 32'b010001_00000_01000_0000000000000110; // m[r[0] + 6] = r[8]
		hd[869] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[870] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[871] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[872] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[873] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[874] <= 32'b101000_0000000000_0000000000010100; // lcd_msg = 20
		hd[875] <= 32'b011000_00000_01000_0000000000000000; // r[8] = SWITCHES
		hd[876] <= 32'b010001_00000_01000_0000000010000101; // m[r[0] + 133] = r[8]
		hd[877] <= 32'b001111_00000_01000_0000000010000101; // r[8] = m[r[0] + 133]
		hd[878] <= 32'b000010_01000_11011_0000000000000000; // r[27] = r[8] + 0
		hd[879] <= 32'b011001_11011_000000000000000000000; // LEDS = r[27]
		hd[880] <= 32'b001111_00000_01000_0000000010000101; // r[8] = m[r[0] + 133]
		hd[881] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[882] <= 32'b011011_11110_01000_0000000000000000; // stack[$sp + 0] = r[8]
		hd[883] <= 32'b011010_00000000000000000000101010; // jump to 42(check_ID), $ra = PC + 1
		hd[884] <= 32'b010000_00000_01001_0000000000000001; // r[9] = 1
		hd[885] <= 32'b011111_11101_01001_01010_00000_000000; // (r[29] != r[9]) ? r[10] = 1 : r[10] = 0
		hd[886] <= 32'b010010_00000_01010_0000001101111011; // if(r[0] == r[10]) jump to 891(L67)
		hd[887] <= 32'b101000_0000000000_0000000000010000; // lcd_msg = 16
		hd[888] <= 32'b011000_00000_01001_0000000000000000; // r[9] = SWITCHES
		hd[889] <= 32'b010001_00000_01001_0000000010000101; // m[r[0] + 133] = r[9]
		hd[890] <= 32'b010100_00000000000000001101110000; // jump to 880(L66)
		hd[891] <= 32'b010000_00000_01001_0000000000000001; // r[9] = 1
		hd[892] <= 32'b010001_00000_01001_0000000010000100; // m[r[0] + 132] = r[9]
		hd[893] <= 32'b001111_00000_01001_0000000010000100; // r[9] = m[r[0] + 132]
		hd[894] <= 32'b001111_00000_01010_0000000000000000; // r[10] = m[r[0] + 0]
		hd[895] <= 32'b000110_01001_01010_01011_00000_000000; // (r[9] < r[10]) ? r[11] = 1 : r[11] = 0
		hd[896] <= 32'b010010_00000_01011_0000001110011110; // if(r[0] == r[11]) jump to 926(L70)
		hd[897] <= 32'b010000_00000_01001_0000000000000111; // r[9] = 7
		hd[898] <= 32'b001111_00000_01010_0000000010000100; // r[10] = m[r[0] + 132]
		hd[899] <= 32'b000000_01001_01010_01001_00000_000000; // r[9] = r[9] + r[10]
		hd[900] <= 32'b001111_01001_01010_0000000000000000; // r[10] = m[r[9] + 0]
		hd[901] <= 32'b001111_00000_01001_0000000010000101; // r[9] = m[r[0] + 133]
		hd[902] <= 32'b011110_01010_01001_01100_00000_000000; // (r[10] == r[9]) ? r[12] = 1 : r[12] = 0
		hd[903] <= 32'b010010_00000_01100_0000001110011010; // if(r[0] == r[12]) jump to 922(L72)
		hd[904] <= 32'b010000_00000_01001_0000000000000111; // r[9] = 7
		hd[905] <= 32'b001111_00000_01010_0000000010000100; // r[10] = m[r[0] + 132]
		hd[906] <= 32'b000000_01001_01010_01001_00000_000000; // r[9] = r[9] + r[10]
		hd[907] <= 32'b010000_00000_01010_0000000001100011; // r[10] = 99
		hd[908] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[909] <= 32'b010000_00000_01001_0000000000010110; // r[9] = 22
		hd[910] <= 32'b001111_00000_01010_0000000010000100; // r[10] = m[r[0] + 132]
		hd[911] <= 32'b000000_01001_01010_01001_00000_000000; // r[9] = r[9] + r[10]
		hd[912] <= 32'b010000_00000_01010_0000000000000000; // r[10] = 0
		hd[913] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[914] <= 32'b010000_00000_01001_0000000000100101; // r[9] = 37
		hd[915] <= 32'b001111_00000_01010_0000000010000100; // r[10] = m[r[0] + 132]
		hd[916] <= 32'b000000_01001_01010_01001_00000_000000; // r[9] = r[9] + r[10]
		hd[917] <= 32'b010000_00000_01010_0000000000000000; // r[10] = 0
		hd[918] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[919] <= 32'b001111_00000_01001_0000000000000000; // r[9] = m[r[0] + 0]
		hd[920] <= 32'b010001_00000_01001_0000000010000100; // m[r[0] + 132] = r[9]
		hd[921] <= 32'b010100_00000000000000001110011101; // jump to 925(L73)
		hd[922] <= 32'b001111_00000_01001_0000000010000100; // r[9] = m[r[0] + 132]
		hd[923] <= 32'b000010_01001_01001_0000000000000001; // r[9] = r[9] + 1
		hd[924] <= 32'b010001_00000_01001_0000000010000100; // m[r[0] + 132] = r[9]
		hd[925] <= 32'b010100_00000000000000001101111101; // jump to 893(L69)
		hd[926] <= 32'b101000_0000000000_0000000000010101; // lcd_msg = 21
		hd[927] <= 32'b011000_00000_01001_0000000000000000; // r[9] = SWITCHES
		hd[928] <= 32'b010001_00000_01001_0000000000000110; // m[r[0] + 6] = r[9]
		hd[929] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[930] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[931] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[932] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[933] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[934] <= 32'b101000_0000000000_0000000000000110; // lcd_msg = 6
		hd[935] <= 32'b011000_00000_01001_0000000000000000; // r[9] = SWITCHES
		hd[936] <= 32'b010001_00000_01001_0000000000000110; // m[r[0] + 6] = r[9]
		hd[937] <= 32'b101000_0000000000_0000000000000111; // lcd_msg = 7
		hd[938] <= 32'b011000_00000_01001_0000000000000000; // r[9] = SWITCHES
		hd[939] <= 32'b010001_00000_01001_0000000010001001; // m[r[0] + 137] = r[9]
		hd[940] <= 32'b001111_00000_01001_0000000010001001; // r[9] = m[r[0] + 137]
		hd[941] <= 32'b000010_01001_11011_0000000000000000; // r[27] = r[9] + 0
		hd[942] <= 32'b011001_11011_000000000000000000000; // LEDS = r[27]
		hd[943] <= 32'b001111_00000_01001_0000000010001001; // r[9] = m[r[0] + 137]
		hd[944] <= 32'b010000_00000_01010_0000000000000001; // r[10] = 1
		hd[945] <= 32'b011110_01001_01010_01011_00000_000000; // (r[9] == r[10]) ? r[11] = 1 : r[11] = 0
		hd[946] <= 32'b010010_00000_01011_0000001111000100; // if(r[0] == r[11]) jump to 964(L74)
		hd[947] <= 32'b001111_00000_01001_0000000000000001; // r[9] = m[r[0] + 1]
		hd[948] <= 32'b001111_00000_01010_0000000000000010; // r[10] = m[r[0] + 2]
		hd[949] <= 32'b011110_01001_01010_01100_00000_000000; // (r[9] == r[10]) ? r[12] = 1 : r[12] = 0
		hd[950] <= 32'b010010_00000_01100_0000001110111011; // if(r[0] == r[12]) jump to 955(L75)
		hd[951] <= 32'b101000_0000000000_0000000000001000; // lcd_msg = 8
		hd[952] <= 32'b011000_00000_01001_0000000000000000; // r[9] = SWITCHES
		hd[953] <= 32'b010001_00000_01001_0000000000000110; // m[r[0] + 6] = r[9]
		hd[954] <= 32'b010100_00000000000000001111000100; // jump to 964(L76)
		hd[955] <= 32'b011010_00000000000000001010111110; // jump to 702(get_free_file_position), $ra = PC + 1
		hd[956] <= 32'b010001_00000_11101_0000000010000110; // m[r[0] + 134] = r[29]
		hd[957] <= 32'b001111_00000_01001_0000000010000110; // r[9] = m[r[0] + 134]
		hd[958] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[959] <= 32'b011011_11110_01001_0000000000000000; // stack[$sp + 0] = r[9]
		hd[960] <= 32'b011010_00000000000000001011011100; // jump to 732(create_file), $ra = PC + 1
		hd[961] <= 32'b001111_00000_01001_0000000000000010; // r[9] = m[r[0] + 2]
		hd[962] <= 32'b000010_01001_01001_0000000000000001; // r[9] = r[9] + 1
		hd[963] <= 32'b010001_00000_01001_0000000000000010; // m[r[0] + 2] = r[9]
		hd[964] <= 32'b001111_00000_01001_0000000010001001; // r[9] = m[r[0] + 137]
		hd[965] <= 32'b010000_00000_01010_0000000000000010; // r[10] = 2
		hd[966] <= 32'b011110_01001_01010_01011_00000_000000; // (r[9] == r[10]) ? r[11] = 1 : r[11] = 0
		hd[967] <= 32'b010010_00000_01011_0000001111001001; // if(r[0] == r[11]) jump to 969(L78)
		hd[968] <= 32'b011010_00000000000000001100100101; // jump to 805(rename_file), $ra = PC + 1
		hd[969] <= 32'b001111_00000_01001_0000000010001001; // r[9] = m[r[0] + 137]
		hd[970] <= 32'b010000_00000_01010_0000000000000011; // r[10] = 3
		hd[971] <= 32'b011110_01001_01010_01011_00000_000000; // (r[9] == r[10]) ? r[11] = 1 : r[11] = 0
		hd[972] <= 32'b010010_00000_01011_0000001111010001; // if(r[0] == r[11]) jump to 977(L80)
		hd[973] <= 32'b011010_00000000000000001101101000; // jump to 872(delete_file), $ra = PC + 1
		hd[974] <= 32'b001111_00000_01001_0000000000000010; // r[9] = m[r[0] + 2]
		hd[975] <= 32'b000011_01001_01001_0000000000000001; // r[9] = r[9] - 1
		hd[976] <= 32'b010001_00000_01001_0000000000000010; // m[r[0] + 2] = r[9]
		hd[977] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[978] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[979] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[980] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[981] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[982] <= 32'b101000_0000000000_0000000000000001; // lcd_msg = 1
		hd[983] <= 32'b011000_00000_01001_0000000000000000; // r[9] = SWITCHES
		hd[984] <= 32'b010001_00000_01001_0000000010001010; // m[r[0] + 138] = r[9]
		hd[985] <= 32'b001111_00000_01001_0000000010001010; // r[9] = m[r[0] + 138]
		hd[986] <= 32'b000010_01001_11011_0000000000000000; // r[27] = r[9] + 0
		hd[987] <= 32'b011001_11011_000000000000000000000; // LEDS = r[27]
		hd[988] <= 32'b001111_00000_01001_0000000010001010; // r[9] = m[r[0] + 138]
		hd[989] <= 32'b010000_00000_01010_0000000000000001; // r[10] = 1
		hd[990] <= 32'b011110_01001_01010_01011_00000_000000; // (r[9] == r[10]) ? r[11] = 1 : r[11] = 0
		hd[991] <= 32'b010010_00000_01011_0000001111100001; // if(r[0] == r[11]) jump to 993(L82)
		hd[992] <= 32'b011010_00000000000000001010001000; // jump to 648(process_operation), $ra = PC + 1
		hd[993] <= 32'b001111_00000_01001_0000000010001010; // r[9] = m[r[0] + 138]
		hd[994] <= 32'b010000_00000_01010_0000000000000010; // r[10] = 2
		hd[995] <= 32'b011110_01001_01010_01011_00000_000000; // (r[9] == r[10]) ? r[11] = 1 : r[11] = 0
		hd[996] <= 32'b010010_00000_01011_0000001111100110; // if(r[0] == r[11]) jump to 998(L84)
		hd[997] <= 32'b011010_00000000000000001110100100; // jump to 932(file_operation), $ra = PC + 1
		hd[998] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[999] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[1000] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[1001] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[1002] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[1003] <= 32'b010000_00000_01001_0000000000001111; // r[9] = 15
		hd[1004] <= 32'b010001_00000_01001_0000000000000000; // m[r[0] + 0] = r[9]
		hd[1005] <= 32'b010000_00000_01001_0000000000001111; // r[9] = 15
		hd[1006] <= 32'b010001_00000_01001_0000000000000001; // m[r[0] + 1] = r[9]
		hd[1007] <= 32'b010000_00000_01001_0000000000001010; // r[9] = 10
		hd[1008] <= 32'b010001_00000_01001_0000000000000010; // m[r[0] + 2] = r[9]
		hd[1009] <= 32'b010000_00000_01001_0000010000000000; // r[9] = 1024
		hd[1010] <= 32'b010001_00000_01001_0000000000000100; // m[r[0] + 4] = r[9]
		hd[1011] <= 32'b010000_00000_01001_0000000011111100; // r[9] = 252
		hd[1012] <= 32'b010001_00000_01001_0000000000000101; // m[r[0] + 5] = r[9]
		hd[1013] <= 32'b010000_00000_01001_0000000000000001; // r[9] = 1
		hd[1014] <= 32'b010001_00000_01001_0000000010001011; // m[r[0] + 139] = r[9]
		hd[1015] <= 32'b001111_00000_01001_0000000010001011; // r[9] = m[r[0] + 139]
		hd[1016] <= 32'b001111_00000_01010_0000000000000000; // r[10] = m[r[0] + 0]
		hd[1017] <= 32'b000110_01001_01010_01011_00000_000000; // (r[9] < r[10]) ? r[11] = 1 : r[11] = 0
		hd[1018] <= 32'b010010_00000_01011_0000010000010011; // if(r[0] == r[11]) jump to 1043(L87)
		hd[1019] <= 32'b001111_00000_01001_0000000010001011; // r[9] = m[r[0] + 139]
		hd[1020] <= 32'b010000_00000_01010_0000000000001010; // r[10] = 10
		hd[1021] <= 32'b000110_01001_01010_01100_00000_000000; // (r[9] < r[10]) ? r[12] = 1 : r[12] = 0
		hd[1022] <= 32'b010010_00000_01100_0000010000000101; // if(r[0] == r[12]) jump to 1029(L89)
		hd[1023] <= 32'b010000_00000_01001_0000000000000111; // r[9] = 7
		hd[1024] <= 32'b001111_00000_01010_0000000010001011; // r[10] = m[r[0] + 139]
		hd[1025] <= 32'b000000_01001_01010_01001_00000_000000; // r[9] = r[9] + r[10]
		hd[1026] <= 32'b001111_00000_01010_0000000010001011; // r[10] = m[r[0] + 139]
		hd[1027] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[1028] <= 32'b010100_00000000000000010000001010; // jump to 1034(L90)
		hd[1029] <= 32'b010000_00000_01001_0000000000000111; // r[9] = 7
		hd[1030] <= 32'b001111_00000_01010_0000000010001011; // r[10] = m[r[0] + 139]
		hd[1031] <= 32'b000000_01001_01010_01001_00000_000000; // r[9] = r[9] + r[10]
		hd[1032] <= 32'b010000_00000_01010_0000000001100011; // r[10] = 99
		hd[1033] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[1034] <= 32'b010000_00000_01001_0000000001010010; // r[9] = 82
		hd[1035] <= 32'b001111_00000_01010_0000000010001011; // r[10] = m[r[0] + 139]
		hd[1036] <= 32'b000000_01001_01010_01001_00000_000000; // r[9] = r[9] + r[10]
		hd[1037] <= 32'b010000_00000_01010_0000000000000000; // r[10] = 0
		hd[1038] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[1039] <= 32'b001111_00000_01001_0000000010001011; // r[9] = m[r[0] + 139]
		hd[1040] <= 32'b000010_01001_01001_0000000000000001; // r[9] = r[9] + 1
		hd[1041] <= 32'b010001_00000_01001_0000000010001011; // m[r[0] + 139] = r[9]
		hd[1042] <= 32'b010100_00000000000000001111110111; // jump to 1015(L86)
		hd[1043] <= 32'b010000_00000_01001_0000000000010110; // r[9] = 22
		hd[1044] <= 32'b000010_01001_01001_0000000000000000; // r[9] = r[9] + 0
		hd[1045] <= 32'b010000_00000_01010_0000000000000000; // r[10] = 0
		hd[1046] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[1047] <= 32'b010000_00000_01001_0000000000100101; // r[9] = 37
		hd[1048] <= 32'b000010_01001_01001_0000000000000000; // r[9] = r[9] + 0
		hd[1049] <= 32'b010000_00000_01010_0000000000000000; // r[10] = 0
		hd[1050] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[1051] <= 32'b010000_00000_01001_0000000000010110; // r[9] = 22
		hd[1052] <= 32'b000010_01001_01001_0000000000000001; // r[9] = r[9] + 1
		hd[1053] <= 32'b010000_00000_01010_0000000000000000; // r[10] = 0
		hd[1054] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[1055] <= 32'b010000_00000_01001_0000000000100101; // r[9] = 37
		hd[1056] <= 32'b000010_01001_01001_0000000000000001; // r[9] = r[9] + 1
		hd[1057] <= 32'b010000_00000_01010_0000000000110011; // r[10] = 51
		hd[1058] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[1059] <= 32'b010000_00000_01001_0000000000010110; // r[9] = 22
		hd[1060] <= 32'b000010_01001_01001_0000000000000010; // r[9] = r[9] + 2
		hd[1061] <= 32'b010000_00000_01010_0000000000000000; // r[10] = 0
		hd[1062] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[1063] <= 32'b010000_00000_01001_0000000000100101; // r[9] = 37
		hd[1064] <= 32'b000010_01001_01001_0000000000000010; // r[9] = r[9] + 2
		hd[1065] <= 32'b010000_00000_01010_0000000001000100; // r[10] = 68
		hd[1066] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[1067] <= 32'b010000_00000_01001_0000000000010110; // r[9] = 22
		hd[1068] <= 32'b000010_01001_01001_0000000000000011; // r[9] = r[9] + 3
		hd[1069] <= 32'b010000_00000_01010_0000000000000000; // r[10] = 0
		hd[1070] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[1071] <= 32'b010000_00000_01001_0000000000100101; // r[9] = 37
		hd[1072] <= 32'b000010_01001_01001_0000000000000011; // r[9] = r[9] + 3
		hd[1073] <= 32'b010000_00000_01010_0000000001001011; // r[10] = 75
		hd[1074] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[1075] <= 32'b010000_00000_01001_0000000000010110; // r[9] = 22
		hd[1076] <= 32'b000010_01001_01001_0000000000000100; // r[9] = r[9] + 4
		hd[1077] <= 32'b010000_00000_01010_0000000000000000; // r[10] = 0
		hd[1078] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[1079] <= 32'b010000_00000_01001_0000000000100101; // r[9] = 37
		hd[1080] <= 32'b000010_01001_01001_0000000000000100; // r[9] = r[9] + 4
		hd[1081] <= 32'b010000_00000_01010_0000000001001100; // r[10] = 76
		hd[1082] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[1083] <= 32'b010000_00000_01001_0000000000010110; // r[9] = 22
		hd[1084] <= 32'b000010_01001_01001_0000000000000101; // r[9] = r[9] + 5
		hd[1085] <= 32'b010000_00000_01010_0000000000000000; // r[10] = 0
		hd[1086] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[1087] <= 32'b010000_00000_01001_0000000000100101; // r[9] = 37
		hd[1088] <= 32'b000010_01001_01001_0000000000000101; // r[9] = r[9] + 5
		hd[1089] <= 32'b010000_00000_01010_0000000010011010; // r[10] = 154
		hd[1090] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[1091] <= 32'b010000_00000_01001_0000000000010110; // r[9] = 22
		hd[1092] <= 32'b000010_01001_01001_0000000000000110; // r[9] = r[9] + 6
		hd[1093] <= 32'b010000_00000_01010_0000000000000000; // r[10] = 0
		hd[1094] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[1095] <= 32'b010000_00000_01001_0000000000100101; // r[9] = 37
		hd[1096] <= 32'b000010_01001_01001_0000000000000110; // r[9] = r[9] + 6
		hd[1097] <= 32'b010000_00000_01010_0000000001001000; // r[10] = 72
		hd[1098] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[1099] <= 32'b010000_00000_01001_0000000000010110; // r[9] = 22
		hd[1100] <= 32'b000010_01001_01001_0000000000000111; // r[9] = r[9] + 7
		hd[1101] <= 32'b010000_00000_01010_0000000000000000; // r[10] = 0
		hd[1102] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[1103] <= 32'b010000_00000_01001_0000000000100101; // r[9] = 37
		hd[1104] <= 32'b000010_01001_01001_0000000000000111; // r[9] = r[9] + 7
		hd[1105] <= 32'b010000_00000_01010_0000000000000000; // r[10] = 0
		hd[1106] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[1107] <= 32'b010000_00000_01001_0000000000010110; // r[9] = 22
		hd[1108] <= 32'b000010_01001_01001_0000000000001000; // r[9] = r[9] + 8
		hd[1109] <= 32'b010000_00000_01010_0000000000000000; // r[10] = 0
		hd[1110] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[1111] <= 32'b010000_00000_01001_0000000000100101; // r[9] = 37
		hd[1112] <= 32'b000010_01001_01001_0000000000001000; // r[9] = r[9] + 8
		hd[1113] <= 32'b010000_00000_01010_0000000000000000; // r[10] = 0
		hd[1114] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[1115] <= 32'b010000_00000_01001_0000000000010110; // r[9] = 22
		hd[1116] <= 32'b000010_01001_01001_0000000000001001; // r[9] = r[9] + 9
		hd[1117] <= 32'b010000_00000_01010_0000000000000000; // r[10] = 0
		hd[1118] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[1119] <= 32'b010000_00000_01001_0000000000100101; // r[9] = 37
		hd[1120] <= 32'b000010_01001_01001_0000000000001001; // r[9] = r[9] + 9
		hd[1121] <= 32'b010000_00000_01010_0000000000000000; // r[10] = 0
		hd[1122] <= 32'b010001_01001_01010_0000000000000000; // m[r[9] + 0] = r[10]
		hd[1123] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[1124] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[1125] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[1126] <= 32'b011010_00000000000000001111101001; // jump to 1001(init), $ra = PC + 1
		hd[1127] <= 32'b101000_0000000000_0000000000000000; // lcd_msg = 0
		hd[1128] <= 32'b011000_00000_01001_0000000000000000; // r[9] = SWITCHES
		hd[1129] <= 32'b010001_00000_01001_0000000000000110; // m[r[0] + 6] = r[9]
		hd[1130] <= 32'b010000_00000_01001_0000000000000001; // r[9] = 1
		hd[1131] <= 32'b001111_00000_01010_0000000000000000; // r[10] = m[r[0] + 0]
		hd[1132] <= 32'b000110_01001_01010_01011_00000_000000; // (r[9] < r[10]) ? r[11] = 1 : r[11] = 0
		hd[1133] <= 32'b010010_00000_01011_0000010001110000; // if(r[0] == r[11]) jump to 1136(L92)
		hd[1134] <= 32'b011010_00000000000000001111010100; // jump to 980(bash), $ra = PC + 1
		hd[1135] <= 32'b010100_00000000000000010001101010; // jump to 1130(L91)
		hd[1136] <= 32'b010110_00000000000000000000000000; // nop
		hd[1137] <= 32'b111111_00000000000000000000000000; // end of the program
		hd[1138] <= 32'b010110_00000000000000000000000000; // nop
		hd[1139] <= 32'b010111_11111111111111111111111111; // hlt




		//prog 1 - pow: stack = 100, mem_loc = 283(252+32-1)- ok
		/*
		hd[2048] <= 32'b010000_00000_11110_0000000001100100; // $sp = 100
		hd[2049] <= 32'b010100_00000000000000000000011110; // jump to 30(main)
		hd[2050] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[2051] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[2052] <= 32'b010001_00000_00001_0000000100011100; // m[r[0] + 284] = r[1]
		hd[2053] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[2054] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[2055] <= 32'b010001_00000_00001_0000000100011011; // m[r[0] + 283] = r[1]
		hd[2056] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[2057] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[2058] <= 32'b010000_00000_00001_0000000000000001; // r[1] = 1
		hd[2059] <= 32'b010001_00000_00001_0000000100011110; // m[r[0] + 286] = r[1]
		hd[2060] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		hd[2061] <= 32'b010001_00000_00001_0000000100011101; // m[r[0] + 285] = r[1]
		hd[2062] <= 32'b001111_00000_00001_0000000100011101; // r[1] = m[r[0] + 285]
		hd[2063] <= 32'b001111_00000_00010_0000000100011100; // r[2] = m[r[0] + 284]
		hd[2064] <= 32'b000110_00001_00010_00011_00000_000000; // (r[1] < r[2]) ? r[3] = 1 : r[3] = 0
		hd[2065] <= 32'b010010_00000_00011_0000000000011010; // if(r[0] == r[3]) jump to 26(L3)
		hd[2066] <= 32'b001111_00000_00001_0000000100011110; // r[1] = m[r[0] + 286]
		hd[2067] <= 32'b001111_00000_00010_0000000100011011; // r[2] = m[r[0] + 283]
		hd[2068] <= 32'b001101_00001_00010_00001_00000_000000; // r[1] = r[1] * r[2]
		hd[2069] <= 32'b010001_00000_00001_0000000100011110; // m[r[0] + 286] = r[1]
		hd[2070] <= 32'b001111_00000_00001_0000000100011101; // r[1] = m[r[0] + 285]
		hd[2071] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[2072] <= 32'b010001_00000_00001_0000000100011101; // m[r[0] + 285] = r[1]
		hd[2073] <= 32'b010100_00000000000000000000001110; // jump to 14(L2)
		hd[2074] <= 32'b001111_00000_11101_0000000100011110; // r[29] = m[r[0] + 286]
		hd[2075] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[2076] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[2077] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[2078] <= 32'b111110_0000000000_0000000000000000; // input syscall
		hd[2079] <= 32'b010110_00000000000000000000000000; // nop
		hd[2080] <= 32'b010001_00000_11011_0000000100011111; // m[r[0] + 287] = r[27]
		hd[2081] <= 32'b111110_0000000000_0000000000000000; // input syscall
		hd[2082] <= 32'b010110_00000000000000000000000000; // nop
		hd[2083] <= 32'b010001_00000_11011_0000000100100000; // m[r[0] + 288] = r[27]
		hd[2084] <= 32'b001111_00000_00001_0000000100011111; // r[1] = m[r[0] + 287]
		hd[2085] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[2086] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[2087] <= 32'b001111_00000_00001_0000000100100000; // r[1] = m[r[0] + 288]
		hd[2088] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[2089] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[2090] <= 32'b011010_00000000000000000000000010; // jump to 2(pow), $ra = PC + 1
		hd[2091] <= 32'b010001_00000_11101_0000000100011111; // m[r[0] + 287] = r[29]
		hd[2092] <= 32'b001111_00000_00001_0000000100011111; // r[1] = m[r[0] + 287]
		hd[2093] <= 32'b000010_00001_11011_0000000000000000; // r[27] = r[1] + 0
		hd[2094] <= 32'b111110_0000000000_0000000000000001; // output syscall
		hd[2095] <= 32'b010110_00000000000000000000000000; // nop
		hd[2096] <= 32'b111111_00000000000000000000000000; // end of the program
		hd[2097] <= 32'b010110_00000000000000000000000000; // nop
		hd[2098] <= 32'b010111_11111111111111111111111111; // hlt
		*/
		
		//prog 1 - pow: stack = 100, mem_loc = 283(252+32-1), NET
		hd[2048] <= 32'b010000_00000_11110_0000000001100100; // $sp = 100
		hd[2049] <= 32'b010100_00000000000000000000011110; // jump to 30(main)
		hd[2050] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[2051] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[2052] <= 32'b010001_00000_00001_0000000100011100; // m[r[0] + 284] = r[1]
		hd[2053] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[2054] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[2055] <= 32'b010001_00000_00001_0000000100011011; // m[r[0] + 283] = r[1]
		hd[2056] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[2057] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[2058] <= 32'b010000_00000_00001_0000000000000001; // r[1] = 1
		hd[2059] <= 32'b010001_00000_00001_0000000100011110; // m[r[0] + 286] = r[1]
		hd[2060] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		hd[2061] <= 32'b010001_00000_00001_0000000100011101; // m[r[0] + 285] = r[1]
		hd[2062] <= 32'b001111_00000_00001_0000000100011101; // r[1] = m[r[0] + 285]
		hd[2063] <= 32'b001111_00000_00010_0000000100011100; // r[2] = m[r[0] + 284]
		hd[2064] <= 32'b000110_00001_00010_00011_00000_000000; // (r[1] < r[2]) ? r[3] = 1 : r[3] = 0
		hd[2065] <= 32'b010010_00000_00011_0000000000011010; // if(r[0] == r[3]) jump to 26(L3)
		hd[2066] <= 32'b001111_00000_00001_0000000100011110; // r[1] = m[r[0] + 286]
		hd[2067] <= 32'b001111_00000_00010_0000000100011011; // r[2] = m[r[0] + 283]
		hd[2068] <= 32'b001101_00001_00010_00001_00000_000000; // r[1] = r[1] * r[2]
		hd[2069] <= 32'b010001_00000_00001_0000000100011110; // m[r[0] + 286] = r[1]
		hd[2070] <= 32'b001111_00000_00001_0000000100011101; // r[1] = m[r[0] + 285]
		hd[2071] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[2072] <= 32'b010001_00000_00001_0000000100011101; // m[r[0] + 285] = r[1]
		hd[2073] <= 32'b010100_00000000000000000000001110; // jump to 14(L2)
		hd[2074] <= 32'b001111_00000_11101_0000000100011110; // r[29] = m[r[0] + 286]
		hd[2075] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[2076] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[2077] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[2078] <= 32'b111110_0000000000_0000000000000010; // uart_input syscall
		hd[2079] <= 32'b010110_00000000000000000000000000; // nop
		hd[2080] <= 32'b010001_00000_11011_0000000100011111; // m[r[0] + 287] = r[27]
		hd[2081] <= 32'b111110_0000000000_0000000000000000; // input syscall
		hd[2082] <= 32'b010110_00000000000000000000000000; // nop
		hd[2083] <= 32'b010001_00000_11011_0000000100100000; // m[r[0] + 288] = r[27]
		hd[2084] <= 32'b001111_00000_00001_0000000100011111; // r[1] = m[r[0] + 287]
		hd[2085] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[2086] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[2087] <= 32'b001111_00000_00001_0000000100100000; // r[1] = m[r[0] + 288]
		hd[2088] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[2089] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[2090] <= 32'b011010_00000000000000000000000010; // jump to 2(pow), $ra = PC + 1
		hd[2091] <= 32'b010001_00000_11101_0000000100011111; // m[r[0] + 287] = r[29]
		hd[2092] <= 32'b001111_00000_00001_0000000100011111; // r[1] = m[r[0] + 287]
		hd[2093] <= 32'b000010_00001_11011_0000000000000000; // r[27] = r[1] + 0
		hd[2094] <= 32'b111110_0000000000_0000000000000011; // uart_output syscall
		hd[2095] <= 32'b010110_00000000000000000000000000; // nop
		hd[2096] <= 32'b010110_00000000000000000000000000; // nop
		hd[2097] <= 32'b111111_00000000000000000000000000; // end of the program
		hd[2098] <= 32'b010110_00000000000000000000000000; // nop
		hd[2099] <= 32'b010111_11111111111111111111111111; // hlt

		//prog 2 - fib: stack = 200, mem_loc = 543(512+32-1)- ok
		/*
		hd[4096] <= 32'b010000_00000_11110_0000000011001000; // $sp = 200
		hd[4097] <= 32'b010100_00000000000000000000101110; // jump to 46(main)
		hd[4098] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[4099] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[4100] <= 32'b010001_00000_00001_0000001000100000; // m[r[0] + 544] = r[1]
		hd[4101] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[4102] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[4103] <= 32'b010001_00000_00001_0000001000011111; // m[r[0] + 543] = r[1]
		hd[4104] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[4105] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[4106] <= 32'b010000_00000_00001_0000000000000010; // r[1] = 2
		hd[4107] <= 32'b010001_00000_00001_0000001000100001; // m[r[0] + 545] = r[1]
		hd[4108] <= 32'b001111_00000_00001_0000001000011111; // r[1] = m[r[0] + 543]
		hd[4109] <= 32'b000010_00001_00001_0000000000000000; // r[1] = r[1] + 0
		hd[4110] <= 32'b010000_00000_00010_0000000000000000; // r[2] = 0
		hd[4111] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[4112] <= 32'b001111_00000_00001_0000001000011111; // r[1] = m[r[0] + 543]
		hd[4113] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[4114] <= 32'b010000_00000_00010_0000000000000001; // r[2] = 1
		hd[4115] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[4116] <= 32'b001111_00000_00001_0000001000100001; // r[1] = m[r[0] + 545]
		hd[4117] <= 32'b001111_00000_00010_0000001000100000; // r[2] = m[r[0] + 544]
		hd[4118] <= 32'b000110_00001_00010_00011_00000_000000; // (r[1] < r[2]) ? r[3] = 1 : r[3] = 0
		hd[4119] <= 32'b010010_00000_00011_0000000000101011; // if(r[0] == r[3]) jump to 43(L3)
		hd[4120] <= 32'b001111_00000_00001_0000001000100001; // r[1] = m[r[0] + 545]
		hd[4121] <= 32'b000011_00001_00001_0000000000000010; // r[1] = r[1] - 2
		hd[4122] <= 32'b001111_00000_00010_0000001000011111; // r[2] = m[r[0] + 543]
		hd[4123] <= 32'b000000_00010_00001_00010_00000_000000; // r[2] = r[2] + r[1]
		hd[4124] <= 32'b001111_00000_00001_0000001000100001; // r[1] = m[r[0] + 545]
		hd[4125] <= 32'b000011_00001_00001_0000000000000001; // r[1] = r[1] - 1
		hd[4126] <= 32'b001111_00000_00100_0000001000011111; // r[4] = m[r[0] + 543]
		hd[4127] <= 32'b000000_00100_00001_00100_00000_000000; // r[4] = r[4] + r[1]
		hd[4128] <= 32'b001111_00100_00001_0000000000000000; // r[1] = m[r[4] + 0]
		hd[4129] <= 32'b001111_00010_00101_0000000000000000; // r[5] = m[r[2] + 0]
		hd[4130] <= 32'b000000_00001_00101_00001_00000_000000; // r[1] = r[1] + r[5]
		hd[4131] <= 32'b001111_00000_00010_0000001000011111; // r[2] = m[r[0] + 543]
		hd[4132] <= 32'b001111_00000_00100_0000001000100001; // r[4] = m[r[0] + 545]
		hd[4133] <= 32'b000000_00010_00100_00010_00000_000000; // r[2] = r[2] + r[4]
		hd[4134] <= 32'b010001_00010_00001_0000000000000000; // m[r[2] + 0] = r[1]
		hd[4135] <= 32'b001111_00000_00001_0000001000100001; // r[1] = m[r[0] + 545]
		hd[4136] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[4137] <= 32'b010001_00000_00001_0000001000100001; // m[r[0] + 545] = r[1]
		hd[4138] <= 32'b010100_00000000000000000000010100; // jump to 20(L2)
		hd[4139] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[4140] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[4141] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[4142] <= 32'b010000_00000_00001_0000000000001010; // r[1] = 10
		hd[4143] <= 32'b010001_00000_00001_0000001000100010; // m[r[0] + 546] = r[1]
		hd[4144] <= 32'b010000_00000_00001_0000001000100100; // r[1] = 548
		hd[4145] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[4146] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[4147] <= 32'b001111_00000_00001_0000001000100010; // r[1] = m[r[0] + 546]
		hd[4148] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[4149] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[4150] <= 32'b011010_00000000000000000000000010; // jump to 2(fib), $ra = PC + 1
		hd[4151] <= 32'b111110_0000000000_0000000000000000; // input syscall
		hd[4152] <= 32'b010110_00000000000000000000000000; // nop
		hd[4153] <= 32'b010001_00000_11011_0000001000100011; // m[r[0] + 547] = r[27]
		hd[4154] <= 32'b010000_00000_00001_0000001000100100; // r[1] = 548
		hd[4155] <= 32'b001111_00000_00010_0000001000100011; // r[2] = m[r[0] + 547]
		hd[4156] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[4157] <= 32'b001111_00001_00010_0000000000000000; // r[2] = m[r[1] + 0]
		hd[4158] <= 32'b000010_00010_11011_0000000000000000; // r[27] = r[2] + 0
		hd[4159] <= 32'b111110_0000000000_0000000000000001; // output syscall
		hd[4160] <= 32'b010110_00000000000000000000000000; // nop
		hd[4161] <= 32'b111111_00000000000000000000000000; // end of the program
		hd[4162] <= 32'b010110_00000000000000000000000000; // nop
		hd[4163] <= 32'b010111_11111111111111111111111111; // hlt
		*/

		//prog 2 - fib: stack = 200, mem_loc = 543(512+32-1), NET
		hd[4096] <= 32'b010000_00000_11110_0000000011001000; // $sp = 200
		hd[4097] <= 32'b010100_00000000000000000000101110; // jump to 46(main)
		hd[4098] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[4099] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[4100] <= 32'b010001_00000_00001_0000001000100000; // m[r[0] + 544] = r[1]
		hd[4101] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[4102] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[4103] <= 32'b010001_00000_00001_0000001000011111; // m[r[0] + 543] = r[1]
		hd[4104] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[4105] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[4106] <= 32'b010000_00000_00001_0000000000000010; // r[1] = 2
		hd[4107] <= 32'b010001_00000_00001_0000001000100001; // m[r[0] + 545] = r[1]
		hd[4108] <= 32'b001111_00000_00001_0000001000011111; // r[1] = m[r[0] + 543]
		hd[4109] <= 32'b000010_00001_00001_0000000000000000; // r[1] = r[1] + 0
		hd[4110] <= 32'b010000_00000_00010_0000000000000000; // r[2] = 0
		hd[4111] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[4112] <= 32'b001111_00000_00001_0000001000011111; // r[1] = m[r[0] + 543]
		hd[4113] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[4114] <= 32'b010000_00000_00010_0000000000000001; // r[2] = 1
		hd[4115] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[4116] <= 32'b001111_00000_00001_0000001000100001; // r[1] = m[r[0] + 545]
		hd[4117] <= 32'b001111_00000_00010_0000001000100000; // r[2] = m[r[0] + 544]
		hd[4118] <= 32'b000110_00001_00010_00011_00000_000000; // (r[1] < r[2]) ? r[3] = 1 : r[3] = 0
		hd[4119] <= 32'b010010_00000_00011_0000000000101011; // if(r[0] == r[3]) jump to 43(L3)
		hd[4120] <= 32'b001111_00000_00001_0000001000100001; // r[1] = m[r[0] + 545]
		hd[4121] <= 32'b000011_00001_00001_0000000000000010; // r[1] = r[1] - 2
		hd[4122] <= 32'b001111_00000_00010_0000001000011111; // r[2] = m[r[0] + 543]
		hd[4123] <= 32'b000000_00010_00001_00010_00000_000000; // r[2] = r[2] + r[1]
		hd[4124] <= 32'b001111_00000_00001_0000001000100001; // r[1] = m[r[0] + 545]
		hd[4125] <= 32'b000011_00001_00001_0000000000000001; // r[1] = r[1] - 1
		hd[4126] <= 32'b001111_00000_00100_0000001000011111; // r[4] = m[r[0] + 543]
		hd[4127] <= 32'b000000_00100_00001_00100_00000_000000; // r[4] = r[4] + r[1]
		hd[4128] <= 32'b001111_00100_00001_0000000000000000; // r[1] = m[r[4] + 0]
		hd[4129] <= 32'b001111_00010_00101_0000000000000000; // r[5] = m[r[2] + 0]
		hd[4130] <= 32'b000000_00001_00101_00001_00000_000000; // r[1] = r[1] + r[5]
		hd[4131] <= 32'b001111_00000_00010_0000001000011111; // r[2] = m[r[0] + 543]
		hd[4132] <= 32'b001111_00000_00100_0000001000100001; // r[4] = m[r[0] + 545]
		hd[4133] <= 32'b000000_00010_00100_00010_00000_000000; // r[2] = r[2] + r[4]
		hd[4134] <= 32'b010001_00010_00001_0000000000000000; // m[r[2] + 0] = r[1]
		hd[4135] <= 32'b001111_00000_00001_0000001000100001; // r[1] = m[r[0] + 545]
		hd[4136] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[4137] <= 32'b010001_00000_00001_0000001000100001; // m[r[0] + 545] = r[1]
		hd[4138] <= 32'b010100_00000000000000000000010100; // jump to 20(L2)
		hd[4139] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[4140] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[4141] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[4142] <= 32'b010000_00000_00001_0000000000001010; // r[1] = 10
		hd[4143] <= 32'b010001_00000_00001_0000001000100010; // m[r[0] + 546] = r[1]
		hd[4144] <= 32'b010000_00000_00001_0000001000100100; // r[1] = 548
		hd[4145] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[4146] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[4147] <= 32'b001111_00000_00001_0000001000100010; // r[1] = m[r[0] + 546]
		hd[4148] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[4149] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[4150] <= 32'b011010_00000000000000000000000010; // jump to 2(fib), $ra = PC + 1
		hd[4151] <= 32'b111110_0000000000_0000000000000010; // uart_input syscall
		hd[4152] <= 32'b010110_00000000000000000000000000; // nop
		hd[4153] <= 32'b010001_00000_11011_0000001000100011; // m[r[0] + 547] = r[27]
		hd[4154] <= 32'b010000_00000_00001_0000001000100100; // r[1] = 548
		hd[4155] <= 32'b001111_00000_00010_0000001000100011; // r[2] = m[r[0] + 547]
		hd[4156] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[4157] <= 32'b001111_00001_00010_0000000000000000; // r[2] = m[r[1] + 0]
		hd[4158] <= 32'b000010_00010_11011_0000000000000000; // r[27] = r[2] + 0
		hd[4159] <= 32'b111110_0000000000_0000000000000011; // uart_output syscall
		hd[4160] <= 32'b010110_00000000000000000000000000; // nop
		hd[4161] <= 32'b010110_00000000000000000000000000; // nop
		hd[4162] <= 32'b111111_00000000000000000000000000; // end of the program
		hd[4163] <= 32'b010110_00000000000000000000000000; // nop
		hd[4164] <= 32'b010111_11111111111111111111111111; // hlt

		//prog 3 - max: stack = 300, mem_loc = 787(756+32-1)
		/*
		hd[6144] <= 32'b010000_00000_11110_0000000100101100; // $sp = 300
		hd[6145] <= 32'b010100_00000000000000000000100110; // jump to 38(main)
		hd[6146] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[6147] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[6148] <= 32'b010001_00000_00001_0000001100010100; // m[r[0] + 788] = r[1]
		hd[6149] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[6150] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[6151] <= 32'b010001_00000_00001_0000001100010011; // m[r[0] + 787] = r[1]
		hd[6152] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[6153] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[6154] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		hd[6155] <= 32'b010001_00000_00001_0000001100010101; // m[r[0] + 789] = r[1]
		hd[6156] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		hd[6157] <= 32'b010001_00000_00001_0000001100010110; // m[r[0] + 790] = r[1]
		hd[6158] <= 32'b001111_00000_00001_0000001100010101; // r[1] = m[r[0] + 789]
		hd[6159] <= 32'b001111_00000_00010_0000001100010100; // r[2] = m[r[0] + 788]
		hd[6160] <= 32'b000110_00001_00010_00011_00000_000000; // (r[1] < r[2]) ? r[3] = 1 : r[3] = 0
		hd[6161] <= 32'b010010_00000_00011_0000000000100010; // if(r[0] == r[3]) jump to 34(L3)
		hd[6162] <= 32'b001111_00000_00001_0000001100010011; // r[1] = m[r[0] + 787]
		hd[6163] <= 32'b001111_00000_00010_0000001100010101; // r[2] = m[r[0] + 789]
		hd[6164] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[6165] <= 32'b001111_00000_00010_0000001100010110; // r[2] = m[r[0] + 790]
		hd[6166] <= 32'b001111_00001_00100_0000000000000000; // r[4] = m[r[1] + 0]
		hd[6167] <= 32'b000110_00010_00100_00001_00000_000000; // (r[2] < r[4]) ? r[1] = 1 : r[1] = 0
		hd[6168] <= 32'b010010_00000_00001_0000000000011110; // if(r[0] == r[1]) jump to 30(L5)
		hd[6169] <= 32'b001111_00000_00010_0000001100010011; // r[2] = m[r[0] + 787]
		hd[6170] <= 32'b001111_00000_00100_0000001100010101; // r[4] = m[r[0] + 789]
		hd[6171] <= 32'b000000_00010_00100_00010_00000_000000; // r[2] = r[2] + r[4]
		hd[6172] <= 32'b001111_00010_00100_0000000000000000; // r[4] = m[r[2] + 0]
		hd[6173] <= 32'b010001_00000_00100_0000001100010110; // m[r[0] + 790] = r[4]
		hd[6174] <= 32'b001111_00000_00001_0000001100010101; // r[1] = m[r[0] + 789]
		hd[6175] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[6176] <= 32'b010001_00000_00001_0000001100010101; // m[r[0] + 789] = r[1]
		hd[6177] <= 32'b010100_00000000000000000000001110; // jump to 14(L2)
		hd[6178] <= 32'b001111_00000_11101_0000001100010110; // r[29] = m[r[0] + 790]
		hd[6179] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[6180] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[6181] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[6182] <= 32'b010000_00000_00001_0000000000000101; // r[1] = 5
		hd[6183] <= 32'b010001_00000_00001_0000001100011100; // m[r[0] + 796] = r[1]
		hd[6184] <= 32'b010000_00000_00001_0000001100010111; // r[1] = 791
		hd[6185] <= 32'b000010_00001_00001_0000000000000000; // r[1] = r[1] + 0
		hd[6186] <= 32'b010000_00000_00010_0000000000001101; // r[2] = 13
		hd[6187] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[6188] <= 32'b010000_00000_00001_0000001100010111; // r[1] = 791
		hd[6189] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[6190] <= 32'b010000_00000_00010_0000000000001001; // r[2] = 9
		hd[6191] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[6192] <= 32'b010000_00000_00001_0000001100010111; // r[1] = 791
		hd[6193] <= 32'b000010_00001_00001_0000000000000010; // r[1] = r[1] + 2
		hd[6194] <= 32'b010000_00000_00010_0000000000111000; // r[2] = 56
		hd[6195] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[6196] <= 32'b010000_00000_00001_0000001100010111; // r[1] = 791
		hd[6197] <= 32'b000010_00001_00001_0000000000000011; // r[1] = r[1] + 3
		hd[6198] <= 32'b010000_00000_00010_0000000000101101; // r[2] = 45
		hd[6199] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[6200] <= 32'b010000_00000_00001_0000001100010111; // r[1] = 791
		hd[6201] <= 32'b000010_00001_00001_0000000000000100; // r[1] = r[1] + 4
		hd[6202] <= 32'b010000_00000_00010_0000000000110011; // r[2] = 51
		hd[6203] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[6204] <= 32'b010000_00000_00001_0000001100010111; // r[1] = 791
		hd[6205] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[6206] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[6207] <= 32'b001111_00000_00001_0000001100011100; // r[1] = m[r[0] + 796]
		hd[6208] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[6209] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[6210] <= 32'b011010_00000000000000000000000010; // jump to 2(max), $ra = PC + 1
		hd[6211] <= 32'b000010_11101_00001_0000000000000000; // r[1] = r[29] + 0
		hd[6212] <= 32'b000010_00001_11011_0000000000000000; // r[27] = r[1] + 0
		hd[6213] <= 32'b111110_0000000000_0000000000000001; // output syscall
		hd[6214] <= 32'b010110_00000000000000000000000000; // nop
		hd[6215] <= 32'b010110_00000000000000000000000000; // nop
		hd[6216] <= 32'b111111_00000000000000000000000000; // end of the program
		hd[6217] <= 32'b010110_00000000000000000000000000; // nop
		hd[6218] <= 32'b010111_11111111111111111111111111; // hlt
		*/
		
		//prog 3 - max: stack = 300, mem_loc = 787(756+32-1), NET
		hd[6144] <= 32'b010000_00000_11110_0000000100101100; // $sp = 300
		hd[6145] <= 32'b010100_00000000000000000000100110; // jump to 38(main)
		hd[6146] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[6147] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[6148] <= 32'b010001_00000_00001_0000001100010100; // m[r[0] + 788] = r[1]
		hd[6149] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[6150] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[6151] <= 32'b010001_00000_00001_0000001100010011; // m[r[0] + 787] = r[1]
		hd[6152] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[6153] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[6154] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		hd[6155] <= 32'b010001_00000_00001_0000001100010101; // m[r[0] + 789] = r[1]
		hd[6156] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		hd[6157] <= 32'b010001_00000_00001_0000001100010110; // m[r[0] + 790] = r[1]
		hd[6158] <= 32'b001111_00000_00001_0000001100010101; // r[1] = m[r[0] + 789]
		hd[6159] <= 32'b001111_00000_00010_0000001100010100; // r[2] = m[r[0] + 788]
		hd[6160] <= 32'b000110_00001_00010_00011_00000_000000; // (r[1] < r[2]) ? r[3] = 1 : r[3] = 0
		hd[6161] <= 32'b010010_00000_00011_0000000000100010; // if(r[0] == r[3]) jump to 34(L3)
		hd[6162] <= 32'b001111_00000_00001_0000001100010011; // r[1] = m[r[0] + 787]
		hd[6163] <= 32'b001111_00000_00010_0000001100010101; // r[2] = m[r[0] + 789]
		hd[6164] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[6165] <= 32'b001111_00000_00010_0000001100010110; // r[2] = m[r[0] + 790]
		hd[6166] <= 32'b001111_00001_00100_0000000000000000; // r[4] = m[r[1] + 0]
		hd[6167] <= 32'b000110_00010_00100_00001_00000_000000; // (r[2] < r[4]) ? r[1] = 1 : r[1] = 0
		hd[6168] <= 32'b010010_00000_00001_0000000000011110; // if(r[0] == r[1]) jump to 30(L5)
		hd[6169] <= 32'b001111_00000_00010_0000001100010011; // r[2] = m[r[0] + 787]
		hd[6170] <= 32'b001111_00000_00100_0000001100010101; // r[4] = m[r[0] + 789]
		hd[6171] <= 32'b000000_00010_00100_00010_00000_000000; // r[2] = r[2] + r[4]
		hd[6172] <= 32'b001111_00010_00100_0000000000000000; // r[4] = m[r[2] + 0]
		hd[6173] <= 32'b010001_00000_00100_0000001100010110; // m[r[0] + 790] = r[4]
		hd[6174] <= 32'b001111_00000_00001_0000001100010101; // r[1] = m[r[0] + 789]
		hd[6175] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[6176] <= 32'b010001_00000_00001_0000001100010101; // m[r[0] + 789] = r[1]
		hd[6177] <= 32'b010100_00000000000000000000001110; // jump to 14(L2)
		hd[6178] <= 32'b001111_00000_11101_0000001100010110; // r[29] = m[r[0] + 790]
		hd[6179] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[6180] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[6181] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[6182] <= 32'b010000_00000_00001_0000000000000101; // r[1] = 5
		hd[6183] <= 32'b010001_00000_00001_0000001100011100; // m[r[0] + 796] = r[1]
		hd[6184] <= 32'b010000_00000_00001_0000001100010111; // r[1] = 791
		hd[6185] <= 32'b000010_00001_00001_0000000000000000; // r[1] = r[1] + 0
		hd[6186] <= 32'b010000_00000_00010_0000000000001101; // r[2] = 13
		hd[6187] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[6188] <= 32'b010000_00000_00001_0000001100010111; // r[1] = 791
		hd[6189] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[6190] <= 32'b010000_00000_00010_0000000000001001; // r[2] = 9
		hd[6191] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[6192] <= 32'b010000_00000_00001_0000001100010111; // r[1] = 791
		hd[6193] <= 32'b000010_00001_00001_0000000000000010; // r[1] = r[1] + 2
		hd[6194] <= 32'b010000_00000_00010_0000000000111000; // r[2] = 56
		hd[6195] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[6196] <= 32'b010000_00000_00001_0000001100010111; // r[1] = 791
		hd[6197] <= 32'b000010_00001_00001_0000000000000011; // r[1] = r[1] + 3
		hd[6198] <= 32'b010000_00000_00010_0000000000101101; // r[2] = 45
		hd[6199] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[6200] <= 32'b010000_00000_00001_0000001100010111; // r[1] = 791
		hd[6201] <= 32'b000010_00001_00001_0000000000000100; // r[1] = r[1] + 4
		hd[6202] <= 32'b010000_00000_00010_0000000000110011; // r[2] = 51
		hd[6203] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[6204] <= 32'b010000_00000_00001_0000001100010111; // r[1] = 791
		hd[6205] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[6206] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[6207] <= 32'b001111_00000_00001_0000001100011100; // r[1] = m[r[0] + 796]
		hd[6208] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[6209] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[6210] <= 32'b011010_00000000000000000000000010; // jump to 2(max), $ra = PC + 1
		hd[6211] <= 32'b000010_11101_00001_0000000000000000; // r[1] = r[29] + 0
		hd[6212] <= 32'b000010_00001_11011_0000000000000000; // r[27] = r[1] + 0
		hd[6213] <= 32'b111110_0000000000_0000000000000011; // uart_output syscall
		hd[6214] <= 32'b010110_00000000000000000000000000; // nop
		hd[6215] <= 32'b010110_00000000000000000000000000; // nop
		hd[6216] <= 32'b111111_00000000000000000000000000; // end of the program
		hd[6217] <= 32'b010110_00000000000000000000000000; // nop
		hd[6218] <= 32'b010111_11111111111111111111111111; // hlt

		
		//prog 4 - min: stack = 400, mem_loc = 1039(1008+32-1)
		hd[8192] <= 32'b010000_00000_11110_0000000110010000; // $sp = 400
		hd[8193] <= 32'b010100_00000000000000000000101001; // jump to 41(main)
		hd[8194] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[8195] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[8196] <= 32'b010001_00000_00001_0000010000010000; // m[r[0] + 1040] = r[1]
		hd[8197] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[8198] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[8199] <= 32'b010001_00000_00001_0000010000001111; // m[r[0] + 1039] = r[1]
		hd[8200] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[8201] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[8202] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		hd[8203] <= 32'b010001_00000_00001_0000010000010001; // m[r[0] + 1041] = r[1]
		hd[8204] <= 32'b001111_00000_00001_0000010000001111; // r[1] = m[r[0] + 1039]
		hd[8205] <= 32'b001111_00000_00010_0000010000010001; // r[2] = m[r[0] + 1041]
		hd[8206] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[8207] <= 32'b001111_00001_00010_0000000000000000; // r[2] = m[r[1] + 0]
		hd[8208] <= 32'b010001_00000_00010_0000010000010010; // m[r[0] + 1042] = r[2]
		hd[8209] <= 32'b001111_00000_00001_0000010000010001; // r[1] = m[r[0] + 1041]
		hd[8210] <= 32'b001111_00000_00010_0000010000010000; // r[2] = m[r[0] + 1040]
		hd[8211] <= 32'b000110_00001_00010_00011_00000_000000; // (r[1] < r[2]) ? r[3] = 1 : r[3] = 0
		hd[8212] <= 32'b010010_00000_00011_0000000000100101; // if(r[0] == r[3]) jump to 37(L3)
		hd[8213] <= 32'b001111_00000_00001_0000010000001111; // r[1] = m[r[0] + 1039]
		hd[8214] <= 32'b001111_00000_00010_0000010000010001; // r[2] = m[r[0] + 1041]
		hd[8215] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[8216] <= 32'b001111_00000_00010_0000010000010010; // r[2] = m[r[0] + 1042]
		hd[8217] <= 32'b001111_00001_00100_0000000000000000; // r[4] = m[r[1] + 0]
		hd[8218] <= 32'b000110_00100_00010_00001_00000_000000; // (r[4] < r[2]) ? r[1] = 1 : r[1] = 0
		hd[8219] <= 32'b010010_00000_00001_0000000000100001; // if(r[0] == r[1]) jump to 33(L5)
		hd[8220] <= 32'b001111_00000_00010_0000010000001111; // r[2] = m[r[0] + 1039]
		hd[8221] <= 32'b001111_00000_00100_0000010000010001; // r[4] = m[r[0] + 1041]
		hd[8222] <= 32'b000000_00010_00100_00010_00000_000000; // r[2] = r[2] + r[4]
		hd[8223] <= 32'b001111_00010_00100_0000000000000000; // r[4] = m[r[2] + 0]
		hd[8224] <= 32'b010001_00000_00100_0000010000010010; // m[r[0] + 1042] = r[4]
		hd[8225] <= 32'b001111_00000_00001_0000010000010001; // r[1] = m[r[0] + 1041]
		hd[8226] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[8227] <= 32'b010001_00000_00001_0000010000010001; // m[r[0] + 1041] = r[1]
		hd[8228] <= 32'b010100_00000000000000000000010001; // jump to 17(L2)
		hd[8229] <= 32'b001111_00000_11101_0000010000010010; // r[29] = m[r[0] + 1042]
		hd[8230] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[8231] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[8232] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[8233] <= 32'b010000_00000_00001_0000000000000100; // r[1] = 4
		hd[8234] <= 32'b010001_00000_00001_0000010000010111; // m[r[0] + 1047] = r[1]
		hd[8235] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		hd[8236] <= 32'b010001_00000_00001_0000010000011000; // m[r[0] + 1048] = r[1]
		hd[8237] <= 32'b010000_00000_00001_0000010000010011; // r[1] = 1043
		hd[8238] <= 32'b000010_00001_00001_0000000000000000; // r[1] = r[1] + 0
		hd[8239] <= 32'b010000_00000_00010_0000000000001101; // r[2] = 13
		hd[8240] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[8241] <= 32'b010000_00000_00001_0000010000010011; // r[1] = 1043
		hd[8242] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[8243] <= 32'b010000_00000_00010_0000000000100001; // r[2] = 33
		hd[8244] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[8245] <= 32'b010000_00000_00001_0000010000010011; // r[1] = 1043
		hd[8246] <= 32'b000010_00001_00001_0000000000000010; // r[1] = r[1] + 2
		hd[8247] <= 32'b010000_00000_00010_0000000000001011; // r[2] = 11
		hd[8248] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[8249] <= 32'b010000_00000_00001_0000010000010011; // r[1] = 1043
		hd[8250] <= 32'b000010_00001_00001_0000000000000011; // r[1] = r[1] + 3
		hd[8251] <= 32'b010000_00000_00010_0000000001001011; // r[2] = 75
		hd[8252] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[8253] <= 32'b010000_00000_00001_0000010000010011; // r[1] = 1043
		hd[8254] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[8255] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[8256] <= 32'b001111_00000_00001_0000010000010111; // r[1] = m[r[0] + 1047]
		hd[8257] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[8258] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[8259] <= 32'b011010_00000000000000000000000010; // jump to 2(min), $ra = PC + 1
		hd[8260] <= 32'b000010_11101_00001_0000000000000000; // r[1] = r[29] + 0
		hd[8261] <= 32'b000010_00001_11011_0000000000000000; // r[27] = r[1] + 0
		hd[8262] <= 32'b111110_0000000000_0000000000000001; // output syscall
		hd[8263] <= 32'b010110_00000000000000000000000000; // nop
		hd[8264] <= 32'b010110_00000000000000000000000000; // nop
		hd[8265] <= 32'b111111_00000000000000000000000000; // end of the program
		hd[8266] <= 32'b010110_00000000000000000000000000; // nop
		hd[8267] <= 32'b010111_11111111111111111111111111; // hlt

		//prog 5 - sort: stack = 500, mem_loc = 1291(1260+32-1)
		hd[10240] <= 32'b010000_00000_11110_0000000111110100; // $sp = 500
		hd[10241] <= 32'b010100_00000000000000000001100111; // jump to 103(main)
		hd[10242] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[10243] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[10244] <= 32'b010001_00000_00001_0000010100001101; // m[r[0] + 1293] = r[1]
		hd[10245] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[10246] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[10247] <= 32'b010001_00000_00001_0000010100001100; // m[r[0] + 1292] = r[1]
		hd[10248] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[10249] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[10250] <= 32'b010001_00000_00001_0000010100001011; // m[r[0] + 1291] = r[1]
		hd[10251] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[10252] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[10253] <= 32'b001111_00000_00001_0000010100001100; // r[1] = m[r[0] + 1292]
		hd[10254] <= 32'b010001_00000_00001_0000010100010000; // m[r[0] + 1296] = r[1]
		hd[10255] <= 32'b001111_00000_00001_0000010100001011; // r[1] = m[r[0] + 1291]
		hd[10256] <= 32'b001111_00000_00010_0000010100001100; // r[2] = m[r[0] + 1292]
		hd[10257] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[10258] <= 32'b001111_00001_00010_0000000000000000; // r[2] = m[r[1] + 0]
		hd[10259] <= 32'b010001_00000_00010_0000010100001111; // m[r[0] + 1295] = r[2]
		hd[10260] <= 32'b001111_00000_00001_0000010100001100; // r[1] = m[r[0] + 1292]
		hd[10261] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[10262] <= 32'b010001_00000_00001_0000010100001110; // m[r[0] + 1294] = r[1]
		hd[10263] <= 32'b001111_00000_00001_0000010100001110; // r[1] = m[r[0] + 1294]
		hd[10264] <= 32'b001111_00000_00010_0000010100001101; // r[2] = m[r[0] + 1293]
		hd[10265] <= 32'b000110_00001_00010_00011_00000_000000; // (r[1] < r[2]) ? r[3] = 1 : r[3] = 0
		hd[10266] <= 32'b010010_00000_00011_0000000000101101; // if(r[0] == r[3]) jump to 45(L3)
		hd[10267] <= 32'b001111_00000_00001_0000010100001011; // r[1] = m[r[0] + 1291]
		hd[10268] <= 32'b001111_00000_00010_0000010100001110; // r[2] = m[r[0] + 1294]
		hd[10269] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[10270] <= 32'b001111_00001_00010_0000000000000000; // r[2] = m[r[1] + 0]
		hd[10271] <= 32'b001111_00000_00001_0000010100001111; // r[1] = m[r[0] + 1295]
		hd[10272] <= 32'b000110_00010_00001_00100_00000_000000; // (r[2] < r[1]) ? r[4] = 1 : r[4] = 0
		hd[10273] <= 32'b010010_00000_00100_0000000000101001; // if(r[0] == r[4]) jump to 41(L5)
		hd[10274] <= 32'b001111_00000_00001_0000010100001011; // r[1] = m[r[0] + 1291]
		hd[10275] <= 32'b001111_00000_00010_0000010100001110; // r[2] = m[r[0] + 1294]
		hd[10276] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[10277] <= 32'b001111_00001_00010_0000000000000000; // r[2] = m[r[1] + 0]
		hd[10278] <= 32'b010001_00000_00010_0000010100001111; // m[r[0] + 1295] = r[2]
		hd[10279] <= 32'b001111_00000_00001_0000010100001110; // r[1] = m[r[0] + 1294]
		hd[10280] <= 32'b010001_00000_00001_0000010100010000; // m[r[0] + 1296] = r[1]
		hd[10281] <= 32'b001111_00000_00001_0000010100001110; // r[1] = m[r[0] + 1294]
		hd[10282] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[10283] <= 32'b010001_00000_00001_0000010100001110; // m[r[0] + 1294] = r[1]
		hd[10284] <= 32'b010100_00000000000000000000010111; // jump to 23(L2)
		hd[10285] <= 32'b001111_00000_11101_0000010100010000; // r[29] = m[r[0] + 1296]
		hd[10286] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[10287] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[10288] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[10289] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[10290] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[10291] <= 32'b010001_00000_00001_0000010100010011; // m[r[0] + 1299] = r[1]
		hd[10292] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[10293] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[10294] <= 32'b010001_00000_00001_0000010100010010; // m[r[0] + 1298] = r[1]
		hd[10295] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[10296] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[10297] <= 32'b010001_00000_00001_0000010100010001; // m[r[0] + 1297] = r[1]
		hd[10298] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[10299] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[10300] <= 32'b001111_00000_00001_0000010100010010; // r[1] = m[r[0] + 1298]
		hd[10301] <= 32'b010001_00000_00001_0000010100010100; // m[r[0] + 1300] = r[1]
		hd[10302] <= 32'b001111_00000_00001_0000010100010011; // r[1] = m[r[0] + 1299]
		hd[10303] <= 32'b000011_00001_00001_0000000000000001; // r[1] = r[1] - 1
		hd[10304] <= 32'b001111_00000_00010_0000010100010100; // r[2] = m[r[0] + 1300]
		hd[10305] <= 32'b000110_00010_00001_00100_00000_000000; // (r[2] < r[1]) ? r[4] = 1 : r[4] = 0
		hd[10306] <= 32'b010010_00000_00100_0000000001100100; // if(r[0] == r[4]) jump to 100(L8)
		hd[10307] <= 32'b001111_00000_00001_0000010100010001; // r[1] = m[r[0] + 1297]
		hd[10308] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[10309] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[10310] <= 32'b001111_00000_00001_0000010100010100; // r[1] = m[r[0] + 1300]
		hd[10311] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[10312] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[10313] <= 32'b001111_00000_00001_0000010100010011; // r[1] = m[r[0] + 1299]
		hd[10314] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[10315] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[10316] <= 32'b011010_00000000000000000000000010; // jump to 2(minloc), $ra = PC + 1
		hd[10317] <= 32'b010001_00000_11101_0000010100010101; // m[r[0] + 1301] = r[29]
		hd[10318] <= 32'b001111_00000_00001_0000010100010001; // r[1] = m[r[0] + 1297]
		hd[10319] <= 32'b001111_00000_00010_0000010100010101; // r[2] = m[r[0] + 1301]
		hd[10320] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[10321] <= 32'b001111_00001_00010_0000000000000000; // r[2] = m[r[1] + 0]
		hd[10322] <= 32'b010001_00000_00010_0000010100010110; // m[r[0] + 1302] = r[2]
		hd[10323] <= 32'b001111_00000_00001_0000010100010001; // r[1] = m[r[0] + 1297]
		hd[10324] <= 32'b001111_00000_00010_0000010100010100; // r[2] = m[r[0] + 1300]
		hd[10325] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[10326] <= 32'b001111_00000_00010_0000010100010001; // r[2] = m[r[0] + 1297]
		hd[10327] <= 32'b001111_00000_00101_0000010100010101; // r[5] = m[r[0] + 1301]
		hd[10328] <= 32'b000000_00010_00101_00010_00000_000000; // r[2] = r[2] + r[5]
		hd[10329] <= 32'b001111_00001_00101_0000000000000000; // r[5] = m[r[1] + 0]
		hd[10330] <= 32'b010001_00010_00101_0000000000000000; // m[r[2] + 0] = r[5]
		hd[10331] <= 32'b001111_00000_00001_0000010100010001; // r[1] = m[r[0] + 1297]
		hd[10332] <= 32'b001111_00000_00010_0000010100010100; // r[2] = m[r[0] + 1300]
		hd[10333] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[10334] <= 32'b001111_00000_00010_0000010100010110; // r[2] = m[r[0] + 1302]
		hd[10335] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[10336] <= 32'b001111_00000_00001_0000010100010100; // r[1] = m[r[0] + 1300]
		hd[10337] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[10338] <= 32'b010001_00000_00001_0000010100010100; // m[r[0] + 1300] = r[1]
		hd[10339] <= 32'b010100_00000000000000000000111110; // jump to 62(L7)
		hd[10340] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[10341] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[10342] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[10343] <= 32'b010000_00000_00001_0000000000000101; // r[1] = 5
		hd[10344] <= 32'b010001_00000_00001_0000010100011100; // m[r[0] + 1308] = r[1]
		hd[10345] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		hd[10346] <= 32'b010001_00000_00001_0000010100011101; // m[r[0] + 1309] = r[1]
		hd[10347] <= 32'b001111_00000_00001_0000010100011101; // r[1] = m[r[0] + 1309]
		hd[10348] <= 32'b001111_00000_00010_0000010100011100; // r[2] = m[r[0] + 1308]
		hd[10349] <= 32'b000110_00001_00010_00100_00000_000000; // (r[1] < r[2]) ? r[4] = 1 : r[4] = 0
		hd[10350] <= 32'b010010_00000_00100_0000000001111011; // if(r[0] == r[4]) jump to 123(L11)
		hd[10351] <= 32'b111110_0000000000_0000000000000000; // input syscall
		hd[10352] <= 32'b010110_00000000000000000000000000; // nop
		hd[10353] <= 32'b010001_00000_11011_0000010100011110; // m[r[0] + 1310] = r[27]
		hd[10354] <= 32'b010000_00000_00001_0000010100010111; // r[1] = 1303
		hd[10355] <= 32'b001111_00000_00010_0000010100011101; // r[2] = m[r[0] + 1309]
		hd[10356] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[10357] <= 32'b001111_00000_00010_0000010100011110; // r[2] = m[r[0] + 1310]
		hd[10358] <= 32'b010001_00001_00010_0000000000000000; // m[r[1] + 0] = r[2]
		hd[10359] <= 32'b001111_00000_00001_0000010100011101; // r[1] = m[r[0] + 1309]
		hd[10360] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[10361] <= 32'b010001_00000_00001_0000010100011101; // m[r[0] + 1309] = r[1]
		hd[10362] <= 32'b010100_00000000000000000001101011; // jump to 107(L10)
		hd[10363] <= 32'b010000_00000_00001_0000010100010111; // r[1] = 1303
		hd[10364] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[10365] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[10366] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		hd[10367] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[10368] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[10369] <= 32'b001111_00000_00001_0000010100011100; // r[1] = m[r[0] + 1308]
		hd[10370] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[10371] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[10372] <= 32'b011010_00000000000000000000110001; // jump to 49(sort), $ra = PC + 1
		hd[10373] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		hd[10374] <= 32'b010001_00000_00001_0000010100011101; // m[r[0] + 1309] = r[1]
		hd[10375] <= 32'b001111_00000_00001_0000010100011101; // r[1] = m[r[0] + 1309]
		hd[10376] <= 32'b001111_00000_00010_0000010100011100; // r[2] = m[r[0] + 1308]
		hd[10377] <= 32'b000110_00001_00010_00100_00000_000000; // (r[1] < r[2]) ? r[4] = 1 : r[4] = 0
		hd[10378] <= 32'b010010_00000_00100_0000000010010110; // if(r[0] == r[4]) jump to 150(L14)
		hd[10379] <= 32'b010000_00000_00001_0000010100010111; // r[1] = 1303
		hd[10380] <= 32'b001111_00000_00010_0000010100011101; // r[2] = m[r[0] + 1309]
		hd[10381] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[10382] <= 32'b001111_00001_00010_0000000000000000; // r[2] = m[r[1] + 0]
		hd[10383] <= 32'b000010_00010_11011_0000000000000000; // r[27] = r[2] + 0
		hd[10384] <= 32'b111110_0000000000_0000000000000001; // output syscall
		hd[10385] <= 32'b010110_00000000000000000000000000; // nop
		hd[10386] <= 32'b001111_00000_00001_0000010100011101; // r[1] = m[r[0] + 1309]
		hd[10387] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[10388] <= 32'b010001_00000_00001_0000010100011101; // m[r[0] + 1309] = r[1]
		hd[10389] <= 32'b010100_00000000000000000010000111; // jump to 135(L13)
		hd[10390] <= 32'b010110_00000000000000000000000000; // nop
		hd[10391] <= 32'b111111_00000000000000000000000000; // end of the program
		hd[10392] <= 32'b010110_00000000000000000000000000; // nop
		hd[10393] <= 32'b010111_11111111111111111111111111; // hlt

		// prog 6 - array average: stack = 600, mem_loc = 1543(1512+32-1)
		hd[12288] <= 32'b010000_00000_11110_0000001001011000; // $sp = 600
		hd[12289] <= 32'b010100_00000000000000000000100101; // jump to 37(main)
		hd[12290] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[12291] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[12292] <= 32'b010001_00000_00001_0000011000001000; // m[r[0] + 1544] = r[1]
		hd[12293] <= 32'b011100_11110_00001_0000000000000000; // r[1] = stack[$sp + 0]
		hd[12294] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[12295] <= 32'b010001_00000_00001_0000011000000111; // m[r[0] + 1543] = r[1]
		hd[12296] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[12297] <= 32'b011011_11110_11111_0000000000000000; // stack[$sp + 0] = $ra
		hd[12298] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		hd[12299] <= 32'b010001_00000_00001_0000011000001010; // m[r[0] + 1546] = r[1]
		hd[12300] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		hd[12301] <= 32'b010001_00000_00001_0000011000001001; // m[r[0] + 1545] = r[1]
		hd[12302] <= 32'b001111_00000_00001_0000011000001001; // r[1] = m[r[0] + 1545]
		hd[12303] <= 32'b001111_00000_00010_0000011000001000; // r[2] = m[r[0] + 1544]
		hd[12304] <= 32'b000110_00001_00010_00011_00000_000000; // (r[1] < r[2]) ? r[3] = 1 : r[3] = 0
		hd[12305] <= 32'b010010_00000_00011_0000000000011101; // if(r[0] == r[3]) jump to 29(L3)
		hd[12306] <= 32'b001111_00000_00001_0000011000000111; // r[1] = m[r[0] + 1543]
		hd[12307] <= 32'b001111_00000_00010_0000011000001001; // r[2] = m[r[0] + 1545]
		hd[12308] <= 32'b000000_00001_00010_00001_00000_000000; // r[1] = r[1] + r[2]
		hd[12309] <= 32'b001111_00000_00010_0000011000001010; // r[2] = m[r[0] + 1546]
		hd[12310] <= 32'b001111_00001_00100_0000000000000000; // r[4] = m[r[1] + 0]
		hd[12311] <= 32'b000000_00010_00100_00010_00000_000000; // r[2] = r[2] + r[4]
		hd[12312] <= 32'b010001_00000_00010_0000011000001010; // m[r[0] + 1546] = r[2]
		hd[12313] <= 32'b001111_00000_00001_0000011000001001; // r[1] = m[r[0] + 1545]
		hd[12314] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[12315] <= 32'b010001_00000_00001_0000011000001001; // m[r[0] + 1545] = r[1]
		hd[12316] <= 32'b010100_00000000000000000000001110; // jump to 14(L2)
		hd[12317] <= 32'b001111_00000_00001_0000011000001010; // r[1] = m[r[0] + 1546]
		hd[12318] <= 32'b001111_00000_00010_0000011000001000; // r[2] = m[r[0] + 1544]
		hd[12319] <= 32'b001110_00001_00010_00001_00000_000000; // r[1] = r[1] / r[2]
		hd[12320] <= 32'b010001_00000_00001_0000011000001010; // m[r[0] + 1546] = r[1]
		hd[12321] <= 32'b001111_00000_11101_0000011000001010; // r[29] = m[r[0] + 1546]
		hd[12322] <= 32'b011100_11110_11111_0000000000000000; // $ra = stack[$sp + 0]
		hd[12323] <= 32'b000101_11110_11110_00000_00000_000000; // $sp -= 1
		hd[12324] <= 32'b010101_11111_00000_0000000000000000; // jump to $ra
		hd[12325] <= 32'b010000_00000_00001_0000000000000101; // r[1] = 5
		hd[12326] <= 32'b010001_00000_00001_0000011000010000; // m[r[0] + 1552] = r[1]
		hd[12327] <= 32'b010000_00000_00001_0000000000000000; // r[1] = 0
		hd[12328] <= 32'b010001_00000_00001_0000011000010001; // m[r[0] + 1553] = r[1]
		hd[12329] <= 32'b001111_00000_00001_0000011000010001; // r[1] = m[r[0] + 1553]
		hd[12330] <= 32'b001111_00000_00010_0000011000010000; // r[2] = m[r[0] + 1552]
		hd[12331] <= 32'b000110_00001_00010_00011_00000_000000; // (r[1] < r[2]) ? r[3] = 1 : r[3] = 0
		hd[12332] <= 32'b010010_00000_00011_0000000000111001; // if(r[0] == r[3]) jump to 57(L6)
		hd[12333] <= 32'b001111_00000_00001_0000011000010001; // r[1] = m[r[0] + 1553]
		hd[12334] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[12335] <= 32'b010000_00000_00010_0000000000001010; // r[2] = 10
		hd[12336] <= 32'b001101_00001_00010_00001_00000_000000; // r[1] = r[1] * r[2]
		hd[12337] <= 32'b010000_00000_00010_0000011000001011; // r[2] = 1547
		hd[12338] <= 32'b001111_00000_00100_0000011000010001; // r[4] = m[r[0] + 1553]
		hd[12339] <= 32'b000000_00010_00100_00010_00000_000000; // r[2] = r[2] + r[4]
		hd[12340] <= 32'b010001_00010_00001_0000000000000000; // m[r[2] + 0] = r[1]
		hd[12341] <= 32'b001111_00000_00001_0000011000010001; // r[1] = m[r[0] + 1553]
		hd[12342] <= 32'b000010_00001_00001_0000000000000001; // r[1] = r[1] + 1
		hd[12343] <= 32'b010001_00000_00001_0000011000010001; // m[r[0] + 1553] = r[1]
		hd[12344] <= 32'b010100_00000000000000000000101001; // jump to 41(L5)
		hd[12345] <= 32'b010000_00000_00001_0000011000001011; // r[1] = 1547
		hd[12346] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[12347] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[12348] <= 32'b001111_00000_00001_0000011000010000; // r[1] = m[r[0] + 1552]
		hd[12349] <= 32'b000100_11110_11110_00000_00000_000000; // $sp += 1
		hd[12350] <= 32'b011011_11110_00001_0000000000000000; // stack[$sp + 0] = r[1]
		hd[12351] <= 32'b011010_00000000000000000000000010; // jump to 2(average), $ra = PC + 1
		hd[12352] <= 32'b000010_11101_00001_0000000000000000; // r[1] = r[29] + 0
		hd[12353] <= 32'b000010_00001_11011_0000000000000000; // r[27] = r[1] + 0
		hd[12354] <= 32'b111110_0000000000_0000000000000001; // output syscall
		hd[12355] <= 32'b010110_00000000000000000000000000; // nop
		hd[12356] <= 32'b010110_00000000000000000000000000; // nop
		hd[12357] <= 32'b111111_00000000000000000000000000; // end of the program
		hd[12358] <= 32'b010110_00000000000000000000000000; // nop
		hd[12359] <= 32'b010111_11111111111111111111111111; // hlt
	
	end
	
	always @ ( posedge clk_write )
	begin
		if( write_flag )
			hd[ REGION * proc_num + track_line ] <= input_data;
	end
	
	always @ ( posedge clk_read )
	begin
		hd_output <= hd[ REGION * proc_num + track_line ];
	end

endmodule 

	